netcdf Ta1 {
dimensions:
	time = 3264 ;
	ycoord = 2 ;
	xcoord = 3 ;
variables:
	double time(time) ;
		time:units = "days since 2009-10-01T00.00" ;
	double ycoord(ycoord) ;
		ycoord:units = "meter" ;
	double xcoord(xcoord) ;
		xcoord:units = "meter" ;
	float Ta(xcoord, ycoord, time) ;
		Ta:units = "Degree Celsius" ;
		Ta:missing_value = -9999.f ;
		Ta:long_name = "Air temperature" ;
data:

 time = 0, 0.0416666666666667, 0.0833333333333333, 0.125, 0.166666666666667, 
    0.208333333333333, 0.25, 0.291666666666667, 0.333333333333333, 0.375, 
    0.416666666666667, 0.458333333333333, 0.5, 0.541666666666667, 
    0.583333333333333, 0.625, 0.666666666666667, 0.708333333333333, 0.75, 
    0.791666666666667, 0.833333333333333, 0.875, 0.916666666666667, 
    0.958333333333333, 1, 1.04166666666667, 1.08333333333333, 1.125, 
    1.16666666666667, 1.20833333333333, 1.25, 1.29166666666667, 
    1.33333333333333, 1.375, 1.41666666666667, 1.45833333333333, 1.5, 
    1.54166666666667, 1.58333333333333, 1.625, 1.66666666666667, 
    1.70833333333333, 1.75, 1.79166666666667, 1.83333333333333, 1.875, 
    1.91666666666667, 1.95833333333333, 2, 2.04166666666667, 
    2.08333333333333, 2.125, 2.16666666666667, 2.20833333333333, 2.25, 
    2.29166666666667, 2.33333333333333, 2.375, 2.41666666666667, 
    2.45833333333333, 2.5, 2.54166666666667, 2.58333333333333, 2.625, 
    2.66666666666667, 2.70833333333333, 2.75, 2.79166666666667, 
    2.83333333333333, 2.875, 2.91666666666667, 2.95833333333333, 3, 
    3.04166666666667, 3.08333333333333, 3.125, 3.16666666666667, 
    3.20833333333333, 3.25, 3.29166666666667, 3.33333333333333, 3.375, 
    3.41666666666667, 3.45833333333333, 3.5, 3.54166666666667, 
    3.58333333333333, 3.625, 3.66666666666667, 3.70833333333333, 3.75, 
    3.79166666666667, 3.83333333333333, 3.875, 3.91666666666667, 
    3.95833333333333, 4, 4.04166666666667, 4.08333333333333, 4.125, 
    4.16666666666667, 4.20833333333333, 4.25, 4.29166666666667, 
    4.33333333333333, 4.375, 4.41666666666667, 4.45833333333333, 4.5, 
    4.54166666666667, 4.58333333333333, 4.625, 4.66666666666667, 
    4.70833333333333, 4.75, 4.79166666666667, 4.83333333333333, 4.875, 
    4.91666666666667, 4.95833333333333, 5, 5.04166666666667, 
    5.08333333333333, 5.125, 5.16666666666667, 5.20833333333333, 5.25, 
    5.29166666666667, 5.33333333333333, 5.375, 5.41666666666667, 
    5.45833333333333, 5.5, 5.54166666666667, 5.58333333333333, 5.625, 
    5.66666666666667, 5.70833333333333, 5.75, 5.79166666666667, 
    5.83333333333333, 5.875, 5.91666666666667, 5.95833333333333, 6, 
    6.04166666666667, 6.08333333333333, 6.125, 6.16666666666667, 
    6.20833333333333, 6.25, 6.29166666666667, 6.33333333333333, 6.375, 
    6.41666666666667, 6.45833333333333, 6.5, 6.54166666666667, 
    6.58333333333333, 6.625, 6.66666666666667, 6.70833333333333, 6.75, 
    6.79166666666667, 6.83333333333333, 6.875, 6.91666666666667, 
    6.95833333333333, 7, 7.04166666666667, 7.08333333333333, 7.125, 
    7.16666666666667, 7.20833333333333, 7.25, 7.29166666666667, 
    7.33333333333333, 7.375, 7.41666666666667, 7.45833333333333, 7.5, 
    7.54166666666667, 7.58333333333333, 7.625, 7.66666666666667, 
    7.70833333333333, 7.75, 7.79166666666667, 7.83333333333333, 7.875, 
    7.91666666666667, 7.95833333333333, 8, 8.04166666666667, 
    8.08333333333333, 8.125, 8.16666666666667, 8.20833333333333, 8.25, 
    8.29166666666667, 8.33333333333333, 8.375, 8.41666666666667, 
    8.45833333333333, 8.5, 8.54166666666667, 8.58333333333333, 8.625, 
    8.66666666666667, 8.70833333333333, 8.75, 8.79166666666667, 
    8.83333333333333, 8.875, 8.91666666666667, 8.95833333333333, 9, 
    9.04166666666667, 9.08333333333333, 9.125, 9.16666666666667, 
    9.20833333333333, 9.25, 9.29166666666667, 9.33333333333333, 9.375, 
    9.41666666666667, 9.45833333333333, 9.5, 9.54166666666667, 
    9.58333333333333, 9.625, 9.66666666666667, 9.70833333333333, 9.75, 
    9.79166666666667, 9.83333333333333, 9.875, 9.91666666666667, 
    9.95833333333333, 10, 10.0416666666667, 10.0833333333333, 10.125, 
    10.1666666666667, 10.2083333333333, 10.25, 10.2916666666667, 
    10.3333333333333, 10.375, 10.4166666666667, 10.4583333333333, 10.5, 
    10.5416666666667, 10.5833333333333, 10.625, 10.6666666666667, 
    10.7083333333333, 10.75, 10.7916666666667, 10.8333333333333, 10.875, 
    10.9166666666667, 10.9583333333333, 11, 11.0416666666667, 
    11.0833333333333, 11.125, 11.1666666666667, 11.2083333333333, 11.25, 
    11.2916666666667, 11.3333333333333, 11.375, 11.4166666666667, 
    11.4583333333333, 11.5, 11.5416666666667, 11.5833333333333, 11.625, 
    11.6666666666667, 11.7083333333333, 11.75, 11.7916666666667, 
    11.8333333333333, 11.875, 11.9166666666667, 11.9583333333333, 12, 
    12.0416666666667, 12.0833333333333, 12.125, 12.1666666666667, 
    12.2083333333333, 12.25, 12.2916666666667, 12.3333333333333, 12.375, 
    12.4166666666667, 12.4583333333333, 12.5, 12.5416666666667, 
    12.5833333333333, 12.625, 12.6666666666667, 12.7083333333333, 12.75, 
    12.7916666666667, 12.8333333333333, 12.875, 12.9166666666667, 
    12.9583333333333, 13, 13.0416666666667, 13.0833333333333, 13.125, 
    13.1666666666667, 13.2083333333333, 13.25, 13.2916666666667, 
    13.3333333333333, 13.375, 13.4166666666667, 13.4583333333333, 13.5, 
    13.5416666666667, 13.5833333333333, 13.625, 13.6666666666667, 
    13.7083333333333, 13.75, 13.7916666666667, 13.8333333333333, 13.875, 
    13.9166666666667, 13.9583333333333, 14, 14.0416666666667, 
    14.0833333333333, 14.125, 14.1666666666667, 14.2083333333333, 14.25, 
    14.2916666666667, 14.3333333333333, 14.375, 14.4166666666667, 
    14.4583333333333, 14.5, 14.5416666666667, 14.5833333333333, 14.625, 
    14.6666666666667, 14.7083333333333, 14.75, 14.7916666666667, 
    14.8333333333333, 14.875, 14.9166666666667, 14.9583333333333, 15, 
    15.0416666666667, 15.0833333333333, 15.125, 15.1666666666667, 
    15.2083333333333, 15.25, 15.2916666666667, 15.3333333333333, 15.375, 
    15.4166666666667, 15.4583333333333, 15.5, 15.5416666666667, 
    15.5833333333333, 15.625, 15.6666666666667, 15.7083333333333, 15.75, 
    15.7916666666667, 15.8333333333333, 15.875, 15.9166666666667, 
    15.9583333333333, 16, 16.0416666666667, 16.0833333333333, 16.125, 
    16.1666666666667, 16.2083333333333, 16.25, 16.2916666666667, 
    16.3333333333333, 16.375, 16.4166666666667, 16.4583333333333, 16.5, 
    16.5416666666667, 16.5833333333333, 16.625, 16.6666666666667, 
    16.7083333333333, 16.75, 16.7916666666667, 16.8333333333333, 16.875, 
    16.9166666666667, 16.9583333333333, 17, 17.0416666666667, 
    17.0833333333333, 17.125, 17.1666666666667, 17.2083333333333, 17.25, 
    17.2916666666667, 17.3333333333333, 17.375, 17.4166666666667, 
    17.4583333333333, 17.5, 17.5416666666667, 17.5833333333333, 17.625, 
    17.6666666666667, 17.7083333333333, 17.75, 17.7916666666667, 
    17.8333333333333, 17.875, 17.9166666666667, 17.9583333333333, 18, 
    18.0416666666667, 18.0833333333333, 18.125, 18.1666666666667, 
    18.2083333333333, 18.25, 18.2916666666667, 18.3333333333333, 18.375, 
    18.4166666666667, 18.4583333333333, 18.5, 18.5416666666667, 
    18.5833333333333, 18.625, 18.6666666666667, 18.7083333333333, 18.75, 
    18.7916666666667, 18.8333333333333, 18.875, 18.9166666666667, 
    18.9583333333333, 19, 19.0416666666667, 19.0833333333333, 19.125, 
    19.1666666666667, 19.2083333333333, 19.25, 19.2916666666667, 
    19.3333333333333, 19.375, 19.4166666666667, 19.4583333333333, 19.5, 
    19.5416666666667, 19.5833333333333, 19.625, 19.6666666666667, 
    19.7083333333333, 19.75, 19.7916666666667, 19.8333333333333, 19.875, 
    19.9166666666667, 19.9583333333333, 20, 20.0416666666667, 
    20.0833333333333, 20.125, 20.1666666666667, 20.2083333333333, 20.25, 
    20.2916666666667, 20.3333333333333, 20.375, 20.4166666666667, 
    20.4583333333333, 20.5, 20.5416666666667, 20.5833333333333, 20.625, 
    20.6666666666667, 20.7083333333333, 20.75, 20.7916666666667, 
    20.8333333333333, 20.875, 20.9166666666667, 20.9583333333333, 21, 
    21.0416666666667, 21.0833333333333, 21.125, 21.1666666666667, 
    21.2083333333333, 21.25, 21.2916666666667, 21.3333333333333, 21.375, 
    21.4166666666667, 21.4583333333333, 21.5, 21.5416666666667, 
    21.5833333333333, 21.625, 21.6666666666667, 21.7083333333333, 21.75, 
    21.7916666666667, 21.8333333333333, 21.875, 21.9166666666667, 
    21.9583333333333, 22, 22.0416666666667, 22.0833333333333, 22.125, 
    22.1666666666667, 22.2083333333333, 22.25, 22.2916666666667, 
    22.3333333333333, 22.375, 22.4166666666667, 22.4583333333333, 22.5, 
    22.5416666666667, 22.5833333333333, 22.625, 22.6666666666667, 
    22.7083333333333, 22.75, 22.7916666666667, 22.8333333333333, 22.875, 
    22.9166666666667, 22.9583333333333, 23, 23.0416666666667, 
    23.0833333333333, 23.125, 23.1666666666667, 23.2083333333333, 23.25, 
    23.2916666666667, 23.3333333333333, 23.375, 23.4166666666667, 
    23.4583333333333, 23.5, 23.5416666666667, 23.5833333333333, 23.625, 
    23.6666666666667, 23.7083333333333, 23.75, 23.7916666666667, 
    23.8333333333333, 23.875, 23.9166666666667, 23.9583333333333, 24, 
    24.0416666666667, 24.0833333333333, 24.125, 24.1666666666667, 
    24.2083333333333, 24.25, 24.2916666666667, 24.3333333333333, 24.375, 
    24.4166666666667, 24.4583333333333, 24.5, 24.5416666666667, 
    24.5833333333333, 24.625, 24.6666666666667, 24.7083333333333, 24.75, 
    24.7916666666667, 24.8333333333333, 24.875, 24.9166666666667, 
    24.9583333333333, 25, 25.0416666666667, 25.0833333333333, 25.125, 
    25.1666666666667, 25.2083333333333, 25.25, 25.2916666666667, 
    25.3333333333333, 25.375, 25.4166666666667, 25.4583333333333, 25.5, 
    25.5416666666667, 25.5833333333333, 25.625, 25.6666666666667, 
    25.7083333333333, 25.75, 25.7916666666667, 25.8333333333333, 25.875, 
    25.9166666666667, 25.9583333333333, 26, 26.0416666666667, 
    26.0833333333333, 26.125, 26.1666666666667, 26.2083333333333, 26.25, 
    26.2916666666667, 26.3333333333333, 26.375, 26.4166666666667, 
    26.4583333333333, 26.5, 26.5416666666667, 26.5833333333333, 26.625, 
    26.6666666666667, 26.7083333333333, 26.75, 26.7916666666667, 
    26.8333333333333, 26.875, 26.9166666666667, 26.9583333333333, 27, 
    27.0416666666667, 27.0833333333333, 27.125, 27.1666666666667, 
    27.2083333333333, 27.25, 27.2916666666667, 27.3333333333333, 27.375, 
    27.4166666666667, 27.4583333333333, 27.5, 27.5416666666667, 
    27.5833333333333, 27.625, 27.6666666666667, 27.7083333333333, 27.75, 
    27.7916666666667, 27.8333333333333, 27.875, 27.9166666666667, 
    27.9583333333333, 28, 28.0416666666667, 28.0833333333333, 28.125, 
    28.1666666666667, 28.2083333333333, 28.25, 28.2916666666667, 
    28.3333333333333, 28.375, 28.4166666666667, 28.4583333333333, 28.5, 
    28.5416666666667, 28.5833333333333, 28.625, 28.6666666666667, 
    28.7083333333333, 28.75, 28.7916666666667, 28.8333333333333, 28.875, 
    28.9166666666667, 28.9583333333333, 29, 29.0416666666667, 
    29.0833333333333, 29.125, 29.1666666666667, 29.2083333333333, 29.25, 
    29.2916666666667, 29.3333333333333, 29.375, 29.4166666666667, 
    29.4583333333333, 29.5, 29.5416666666667, 29.5833333333333, 29.625, 
    29.6666666666667, 29.7083333333333, 29.75, 29.7916666666667, 
    29.8333333333333, 29.875, 29.9166666666667, 29.9583333333333, 30, 
    30.0416666666667, 30.0833333333333, 30.125, 30.1666666666667, 
    30.2083333333333, 30.25, 30.2916666666667, 30.3333333333333, 30.375, 
    30.4166666666667, 30.4583333333333, 30.5, 30.5416666666667, 
    30.5833333333333, 30.625, 30.6666666666667, 30.7083333333333, 30.75, 
    30.7916666666667, 30.8333333333333, 30.875, 30.9166666666667, 
    30.9583333333333, 31, 31.0416666666667, 31.0833333333333, 31.125, 
    31.1666666666667, 31.2083333333333, 31.25, 31.2916666666667, 
    31.3333333333333, 31.375, 31.4166666666667, 31.4583333333333, 31.5, 
    31.5416666666667, 31.5833333333333, 31.625, 31.6666666666667, 
    31.7083333333333, 31.75, 31.7916666666667, 31.8333333333333, 31.875, 
    31.9166666666667, 31.9583333333333, 32, 32.0416666666667, 
    32.0833333333333, 32.125, 32.1666666666667, 32.2083333333333, 32.25, 
    32.2916666666667, 32.3333333333333, 32.375, 32.4166666666667, 
    32.4583333333333, 32.5, 32.5416666666667, 32.5833333333333, 32.625, 
    32.6666666666667, 32.7083333333333, 32.75, 32.7916666666667, 
    32.8333333333333, 32.875, 32.9166666666667, 32.9583333333333, 33, 
    33.0416666666667, 33.0833333333333, 33.125, 33.1666666666667, 
    33.2083333333333, 33.25, 33.2916666666667, 33.3333333333333, 33.375, 
    33.4166666666667, 33.4583333333333, 33.5, 33.5416666666667, 
    33.5833333333333, 33.625, 33.6666666666667, 33.7083333333333, 33.75, 
    33.7916666666667, 33.8333333333333, 33.875, 33.9166666666667, 
    33.9583333333333, 34, 34.0416666666667, 34.0833333333333, 34.125, 
    34.1666666666667, 34.2083333333333, 34.25, 34.2916666666667, 
    34.3333333333333, 34.375, 34.4166666666667, 34.4583333333333, 34.5, 
    34.5416666666667, 34.5833333333333, 34.625, 34.6666666666667, 
    34.7083333333333, 34.75, 34.7916666666667, 34.8333333333333, 34.875, 
    34.9166666666667, 34.9583333333333, 35, 35.0416666666667, 
    35.0833333333333, 35.125, 35.1666666666667, 35.2083333333333, 35.25, 
    35.2916666666667, 35.3333333333333, 35.375, 35.4166666666667, 
    35.4583333333333, 35.5, 35.5416666666667, 35.5833333333333, 35.625, 
    35.6666666666667, 35.7083333333333, 35.75, 35.7916666666667, 
    35.8333333333333, 35.875, 35.9166666666667, 35.9583333333333, 36, 
    36.0416666666667, 36.0833333333333, 36.125, 36.1666666666667, 
    36.2083333333333, 36.25, 36.2916666666667, 36.3333333333333, 36.375, 
    36.4166666666667, 36.4583333333333, 36.5, 36.5416666666667, 
    36.5833333333333, 36.625, 36.6666666666667, 36.7083333333333, 36.75, 
    36.7916666666667, 36.8333333333333, 36.875, 36.9166666666667, 
    36.9583333333333, 37, 37.0416666666667, 37.0833333333333, 37.125, 
    37.1666666666667, 37.2083333333333, 37.25, 37.2916666666667, 
    37.3333333333333, 37.375, 37.4166666666667, 37.4583333333333, 37.5, 
    37.5416666666667, 37.5833333333333, 37.625, 37.6666666666667, 
    37.7083333333333, 37.75, 37.7916666666667, 37.8333333333333, 37.875, 
    37.9166666666667, 37.9583333333333, 38, 38.0416666666667, 
    38.0833333333333, 38.125, 38.1666666666667, 38.2083333333333, 38.25, 
    38.2916666666667, 38.3333333333333, 38.375, 38.4166666666667, 
    38.4583333333333, 38.5, 38.5416666666667, 38.5833333333333, 38.625, 
    38.6666666666667, 38.7083333333333, 38.75, 38.7916666666667, 
    38.8333333333333, 38.875, 38.9166666666667, 38.9583333333333, 39, 
    39.0416666666667, 39.0833333333333, 39.125, 39.1666666666667, 
    39.2083333333333, 39.25, 39.2916666666667, 39.3333333333333, 39.375, 
    39.4166666666667, 39.4583333333333, 39.5, 39.5416666666667, 
    39.5833333333333, 39.625, 39.6666666666667, 39.7083333333333, 39.75, 
    39.7916666666667, 39.8333333333333, 39.875, 39.9166666666667, 
    39.9583333333333, 40, 40.0416666666667, 40.0833333333333, 40.125, 
    40.1666666666667, 40.2083333333333, 40.25, 40.2916666666667, 
    40.3333333333333, 40.375, 40.4166666666667, 40.4583333333333, 40.5, 
    40.5416666666667, 40.5833333333333, 40.625, 40.6666666666667, 
    40.7083333333333, 40.75, 40.7916666666667, 40.8333333333333, 40.875, 
    40.9166666666667, 40.9583333333333, 41, 41.0416666666667, 
    41.0833333333333, 41.125, 41.1666666666667, 41.2083333333333, 41.25, 
    41.2916666666667, 41.3333333333333, 41.375, 41.4166666666667, 
    41.4583333333333, 41.5, 41.5416666666667, 41.5833333333333, 41.625, 
    41.6666666666667, 41.7083333333333, 41.75, 41.7916666666667, 
    41.8333333333333, 41.875, 41.9166666666667, 41.9583333333333, 42, 
    42.0416666666667, 42.0833333333333, 42.125, 42.1666666666667, 
    42.2083333333333, 42.25, 42.2916666666667, 42.3333333333333, 42.375, 
    42.4166666666667, 42.4583333333333, 42.5, 42.5416666666667, 
    42.5833333333333, 42.625, 42.6666666666667, 42.7083333333333, 42.75, 
    42.7916666666667, 42.8333333333333, 42.875, 42.9166666666667, 
    42.9583333333333, 43, 43.0416666666667, 43.0833333333333, 43.125, 
    43.1666666666667, 43.2083333333333, 43.25, 43.2916666666667, 
    43.3333333333333, 43.375, 43.4166666666667, 43.4583333333333, 43.5, 
    43.5416666666667, 43.5833333333333, 43.625, 43.6666666666667, 
    43.7083333333333, 43.75, 43.7916666666667, 43.8333333333333, 43.875, 
    43.9166666666667, 43.9583333333333, 44, 44.0416666666667, 
    44.0833333333333, 44.125, 44.1666666666667, 44.2083333333333, 44.25, 
    44.2916666666667, 44.3333333333333, 44.375, 44.4166666666667, 
    44.4583333333333, 44.5, 44.5416666666667, 44.5833333333333, 44.625, 
    44.6666666666667, 44.7083333333333, 44.75, 44.7916666666667, 
    44.8333333333333, 44.875, 44.9166666666667, 44.9583333333333, 45, 
    45.0416666666667, 45.0833333333333, 45.125, 45.1666666666667, 
    45.2083333333333, 45.25, 45.2916666666667, 45.3333333333333, 45.375, 
    45.4166666666667, 45.4583333333333, 45.5, 45.5416666666667, 
    45.5833333333333, 45.625, 45.6666666666667, 45.7083333333333, 45.75, 
    45.7916666666667, 45.8333333333333, 45.875, 45.9166666666667, 
    45.9583333333333, 46, 46.0416666666667, 46.0833333333333, 46.125, 
    46.1666666666667, 46.2083333333333, 46.25, 46.2916666666667, 
    46.3333333333333, 46.375, 46.4166666666667, 46.4583333333333, 46.5, 
    46.5416666666667, 46.5833333333333, 46.625, 46.6666666666667, 
    46.7083333333333, 46.75, 46.7916666666667, 46.8333333333333, 46.875, 
    46.9166666666667, 46.9583333333333, 47, 47.0416666666667, 
    47.0833333333333, 47.125, 47.1666666666667, 47.2083333333333, 47.25, 
    47.2916666666667, 47.3333333333333, 47.375, 47.4166666666667, 
    47.4583333333333, 47.5, 47.5416666666667, 47.5833333333333, 47.625, 
    47.6666666666667, 47.7083333333333, 47.75, 47.7916666666667, 
    47.8333333333333, 47.875, 47.9166666666667, 47.9583333333333, 48, 
    48.0416666666667, 48.0833333333333, 48.125, 48.1666666666667, 
    48.2083333333333, 48.25, 48.2916666666667, 48.3333333333333, 48.375, 
    48.4166666666667, 48.4583333333333, 48.5, 48.5416666666667, 
    48.5833333333333, 48.625, 48.6666666666667, 48.7083333333333, 48.75, 
    48.7916666666667, 48.8333333333333, 48.875, 48.9166666666667, 
    48.9583333333333, 49, 49.0416666666667, 49.0833333333333, 49.125, 
    49.1666666666667, 49.2083333333333, 49.25, 49.2916666666667, 
    49.3333333333333, 49.375, 49.4166666666667, 49.4583333333333, 49.5, 
    49.5416666666667, 49.5833333333333, 49.625, 49.6666666666667, 
    49.7083333333333, 49.75, 49.7916666666667, 49.8333333333333, 49.875, 
    49.9166666666667, 49.9583333333333, 50, 50.0416666666667, 
    50.0833333333333, 50.125, 50.1666666666667, 50.2083333333333, 50.25, 
    50.2916666666667, 50.3333333333333, 50.375, 50.4166666666667, 
    50.4583333333333, 50.5, 50.5416666666667, 50.5833333333333, 50.625, 
    50.6666666666667, 50.7083333333333, 50.75, 50.7916666666667, 
    50.8333333333333, 50.875, 50.9166666666667, 50.9583333333333, 51, 
    51.0416666666667, 51.0833333333333, 51.125, 51.1666666666667, 
    51.2083333333333, 51.25, 51.2916666666667, 51.3333333333333, 51.375, 
    51.4166666666667, 51.4583333333333, 51.5, 51.5416666666667, 
    51.5833333333333, 51.625, 51.6666666666667, 51.7083333333333, 51.75, 
    51.7916666666667, 51.8333333333333, 51.875, 51.9166666666667, 
    51.9583333333333, 52, 52.0416666666667, 52.0833333333333, 52.125, 
    52.1666666666667, 52.2083333333333, 52.25, 52.2916666666667, 
    52.3333333333333, 52.375, 52.4166666666667, 52.4583333333333, 52.5, 
    52.5416666666667, 52.5833333333333, 52.625, 52.6666666666667, 
    52.7083333333333, 52.75, 52.7916666666667, 52.8333333333333, 52.875, 
    52.9166666666667, 52.9583333333333, 53, 53.0416666666667, 
    53.0833333333333, 53.125, 53.1666666666667, 53.2083333333333, 53.25, 
    53.2916666666667, 53.3333333333333, 53.375, 53.4166666666667, 
    53.4583333333333, 53.5, 53.5416666666667, 53.5833333333333, 53.625, 
    53.6666666666667, 53.7083333333333, 53.75, 53.7916666666667, 
    53.8333333333333, 53.875, 53.9166666666667, 53.9583333333333, 54, 
    54.0416666666667, 54.0833333333333, 54.125, 54.1666666666667, 
    54.2083333333333, 54.25, 54.2916666666667, 54.3333333333333, 54.375, 
    54.4166666666667, 54.4583333333333, 54.5, 54.5416666666667, 
    54.5833333333333, 54.625, 54.6666666666667, 54.7083333333333, 54.75, 
    54.7916666666667, 54.8333333333333, 54.875, 54.9166666666667, 
    54.9583333333333, 55, 55.0416666666667, 55.0833333333333, 55.125, 
    55.1666666666667, 55.2083333333333, 55.25, 55.2916666666667, 
    55.3333333333333, 55.375, 55.4166666666667, 55.4583333333333, 55.5, 
    55.5416666666667, 55.5833333333333, 55.625, 55.6666666666667, 
    55.7083333333333, 55.75, 55.7916666666667, 55.8333333333333, 55.875, 
    55.9166666666667, 55.9583333333333, 56, 56.0416666666667, 
    56.0833333333333, 56.125, 56.1666666666667, 56.2083333333333, 56.25, 
    56.2916666666667, 56.3333333333333, 56.375, 56.4166666666667, 
    56.4583333333333, 56.5, 56.5416666666667, 56.5833333333333, 56.625, 
    56.6666666666667, 56.7083333333333, 56.75, 56.7916666666667, 
    56.8333333333333, 56.875, 56.9166666666667, 56.9583333333333, 57, 
    57.0416666666667, 57.0833333333333, 57.125, 57.1666666666667, 
    57.2083333333333, 57.25, 57.2916666666667, 57.3333333333333, 57.375, 
    57.4166666666667, 57.4583333333333, 57.5, 57.5416666666667, 
    57.5833333333333, 57.625, 57.6666666666667, 57.7083333333333, 57.75, 
    57.7916666666667, 57.8333333333333, 57.875, 57.9166666666667, 
    57.9583333333333, 58, 58.0416666666667, 58.0833333333333, 58.125, 
    58.1666666666667, 58.2083333333333, 58.25, 58.2916666666667, 
    58.3333333333333, 58.375, 58.4166666666667, 58.4583333333333, 58.5, 
    58.5416666666667, 58.5833333333333, 58.625, 58.6666666666667, 
    58.7083333333333, 58.75, 58.7916666666667, 58.8333333333333, 58.875, 
    58.9166666666667, 58.9583333333333, 59, 59.0416666666667, 
    59.0833333333333, 59.125, 59.1666666666667, 59.2083333333333, 59.25, 
    59.2916666666667, 59.3333333333333, 59.375, 59.4166666666667, 
    59.4583333333333, 59.5, 59.5416666666667, 59.5833333333333, 59.625, 
    59.6666666666667, 59.7083333333333, 59.75, 59.7916666666667, 
    59.8333333333333, 59.875, 59.9166666666667, 59.9583333333333, 60, 
    60.0416666666667, 60.0833333333333, 60.125, 60.1666666666667, 
    60.2083333333333, 60.25, 60.2916666666667, 60.3333333333333, 60.375, 
    60.4166666666667, 60.4583333333333, 60.5, 60.5416666666667, 
    60.5833333333333, 60.625, 60.6666666666667, 60.7083333333333, 60.75, 
    60.7916666666667, 60.8333333333333, 60.875, 60.9166666666667, 
    60.9583333333333, 61, 61.0416666666667, 61.0833333333333, 61.125, 
    61.1666666666667, 61.2083333333333, 61.25, 61.2916666666667, 
    61.3333333333333, 61.375, 61.4166666666667, 61.4583333333333, 61.5, 
    61.5416666666667, 61.5833333333333, 61.625, 61.6666666666667, 
    61.7083333333333, 61.75, 61.7916666666667, 61.8333333333333, 61.875, 
    61.9166666666667, 61.9583333333333, 62, 62.0416666666667, 
    62.0833333333333, 62.125, 62.1666666666667, 62.2083333333333, 62.25, 
    62.2916666666667, 62.3333333333333, 62.375, 62.4166666666667, 
    62.4583333333333, 62.5, 62.5416666666667, 62.5833333333333, 62.625, 
    62.6666666666667, 62.7083333333333, 62.75, 62.7916666666667, 
    62.8333333333333, 62.875, 62.9166666666667, 62.9583333333333, 63, 
    63.0416666666667, 63.0833333333333, 63.125, 63.1666666666667, 
    63.2083333333333, 63.25, 63.2916666666667, 63.3333333333333, 63.375, 
    63.4166666666667, 63.4583333333333, 63.5, 63.5416666666667, 
    63.5833333333333, 63.625, 63.6666666666667, 63.7083333333333, 63.75, 
    63.7916666666667, 63.8333333333333, 63.875, 63.9166666666667, 
    63.9583333333333, 64, 64.0416666666667, 64.0833333333333, 64.125, 
    64.1666666666667, 64.2083333333333, 64.25, 64.2916666666667, 
    64.3333333333333, 64.375, 64.4166666666667, 64.4583333333333, 64.5, 
    64.5416666666667, 64.5833333333333, 64.625, 64.6666666666667, 
    64.7083333333333, 64.75, 64.7916666666667, 64.8333333333333, 64.875, 
    64.9166666666667, 64.9583333333333, 65, 65.0416666666667, 
    65.0833333333333, 65.125, 65.1666666666667, 65.2083333333333, 65.25, 
    65.2916666666667, 65.3333333333333, 65.375, 65.4166666666667, 
    65.4583333333333, 65.5, 65.5416666666667, 65.5833333333333, 65.625, 
    65.6666666666667, 65.7083333333333, 65.75, 65.7916666666667, 
    65.8333333333333, 65.875, 65.9166666666667, 65.9583333333333, 66, 
    66.0416666666667, 66.0833333333333, 66.125, 66.1666666666667, 
    66.2083333333333, 66.25, 66.2916666666667, 66.3333333333333, 66.375, 
    66.4166666666667, 66.4583333333333, 66.5, 66.5416666666667, 
    66.5833333333333, 66.625, 66.6666666666667, 66.7083333333333, 66.75, 
    66.7916666666667, 66.8333333333333, 66.875, 66.9166666666667, 
    66.9583333333333, 67, 67.0416666666667, 67.0833333333333, 67.125, 
    67.1666666666667, 67.2083333333333, 67.25, 67.2916666666667, 
    67.3333333333333, 67.375, 67.4166666666667, 67.4583333333333, 67.5, 
    67.5416666666667, 67.5833333333333, 67.625, 67.6666666666667, 
    67.7083333333333, 67.75, 67.7916666666667, 67.8333333333333, 67.875, 
    67.9166666666667, 67.9583333333333, 68, 68.0416666666667, 
    68.0833333333333, 68.125, 68.1666666666667, 68.2083333333333, 68.25, 
    68.2916666666667, 68.3333333333333, 68.375, 68.4166666666667, 
    68.4583333333333, 68.5, 68.5416666666667, 68.5833333333333, 68.625, 
    68.6666666666667, 68.7083333333333, 68.75, 68.7916666666667, 
    68.8333333333333, 68.875, 68.9166666666667, 68.9583333333333, 69, 
    69.0416666666667, 69.0833333333333, 69.125, 69.1666666666667, 
    69.2083333333333, 69.25, 69.2916666666667, 69.3333333333333, 69.375, 
    69.4166666666667, 69.4583333333333, 69.5, 69.5416666666667, 
    69.5833333333333, 69.625, 69.6666666666667, 69.7083333333333, 69.75, 
    69.7916666666667, 69.8333333333333, 69.875, 69.9166666666667, 
    69.9583333333333, 70, 70.0416666666667, 70.0833333333333, 70.125, 
    70.1666666666667, 70.2083333333333, 70.25, 70.2916666666667, 
    70.3333333333333, 70.375, 70.4166666666667, 70.4583333333333, 70.5, 
    70.5416666666667, 70.5833333333333, 70.625, 70.6666666666667, 
    70.7083333333333, 70.75, 70.7916666666667, 70.8333333333333, 70.875, 
    70.9166666666667, 70.9583333333333, 71, 71.0416666666667, 
    71.0833333333333, 71.125, 71.1666666666667, 71.2083333333333, 71.25, 
    71.2916666666667, 71.3333333333333, 71.375, 71.4166666666667, 
    71.4583333333333, 71.5, 71.5416666666667, 71.5833333333333, 71.625, 
    71.6666666666667, 71.7083333333333, 71.75, 71.7916666666667, 
    71.8333333333333, 71.875, 71.9166666666667, 71.9583333333333, 72, 
    72.0416666666667, 72.0833333333333, 72.125, 72.1666666666667, 
    72.2083333333333, 72.25, 72.2916666666667, 72.3333333333333, 72.375, 
    72.4166666666667, 72.4583333333333, 72.5, 72.5416666666667, 
    72.5833333333333, 72.625, 72.6666666666667, 72.7083333333333, 72.75, 
    72.7916666666667, 72.8333333333333, 72.875, 72.9166666666667, 
    72.9583333333333, 73, 73.0416666666667, 73.0833333333333, 73.125, 
    73.1666666666667, 73.2083333333333, 73.25, 73.2916666666667, 
    73.3333333333333, 73.375, 73.4166666666667, 73.4583333333333, 73.5, 
    73.5416666666667, 73.5833333333333, 73.625, 73.6666666666667, 
    73.7083333333333, 73.75, 73.7916666666667, 73.8333333333333, 73.875, 
    73.9166666666667, 73.9583333333333, 74, 74.0416666666667, 
    74.0833333333333, 74.125, 74.1666666666667, 74.2083333333333, 74.25, 
    74.2916666666667, 74.3333333333333, 74.375, 74.4166666666667, 
    74.4583333333333, 74.5, 74.5416666666667, 74.5833333333333, 74.625, 
    74.6666666666667, 74.7083333333333, 74.75, 74.7916666666667, 
    74.8333333333333, 74.875, 74.9166666666667, 74.9583333333333, 75, 
    75.0416666666667, 75.0833333333333, 75.125, 75.1666666666667, 
    75.2083333333333, 75.25, 75.2916666666667, 75.3333333333333, 75.375, 
    75.4166666666667, 75.4583333333333, 75.5, 75.5416666666667, 
    75.5833333333333, 75.625, 75.6666666666667, 75.7083333333333, 75.75, 
    75.7916666666667, 75.8333333333333, 75.875, 75.9166666666667, 
    75.9583333333333, 76, 76.0416666666667, 76.0833333333333, 76.125, 
    76.1666666666667, 76.2083333333333, 76.25, 76.2916666666667, 
    76.3333333333333, 76.375, 76.4166666666667, 76.4583333333333, 76.5, 
    76.5416666666667, 76.5833333333333, 76.625, 76.6666666666667, 
    76.7083333333333, 76.75, 76.7916666666667, 76.8333333333333, 76.875, 
    76.9166666666667, 76.9583333333333, 77, 77.0416666666667, 
    77.0833333333333, 77.125, 77.1666666666667, 77.2083333333333, 77.25, 
    77.2916666666667, 77.3333333333333, 77.375, 77.4166666666667, 
    77.4583333333333, 77.5, 77.5416666666667, 77.5833333333333, 77.625, 
    77.6666666666667, 77.7083333333333, 77.75, 77.7916666666667, 
    77.8333333333333, 77.875, 77.9166666666667, 77.9583333333333, 78, 
    78.0416666666667, 78.0833333333333, 78.125, 78.1666666666667, 
    78.2083333333333, 78.25, 78.2916666666667, 78.3333333333333, 78.375, 
    78.4166666666667, 78.4583333333333, 78.5, 78.5416666666667, 
    78.5833333333333, 78.625, 78.6666666666667, 78.7083333333333, 78.75, 
    78.7916666666667, 78.8333333333333, 78.875, 78.9166666666667, 
    78.9583333333333, 79, 79.0416666666667, 79.0833333333333, 79.125, 
    79.1666666666667, 79.2083333333333, 79.25, 79.2916666666667, 
    79.3333333333333, 79.375, 79.4166666666667, 79.4583333333333, 79.5, 
    79.5416666666667, 79.5833333333333, 79.625, 79.6666666666667, 
    79.7083333333333, 79.75, 79.7916666666667, 79.8333333333333, 79.875, 
    79.9166666666667, 79.9583333333333, 80, 80.0416666666667, 
    80.0833333333333, 80.125, 80.1666666666667, 80.2083333333333, 80.25, 
    80.2916666666667, 80.3333333333333, 80.375, 80.4166666666667, 
    80.4583333333333, 80.5, 80.5416666666667, 80.5833333333333, 80.625, 
    80.6666666666667, 80.7083333333333, 80.75, 80.7916666666667, 
    80.8333333333333, 80.875, 80.9166666666667, 80.9583333333333, 81, 
    81.0416666666667, 81.0833333333333, 81.125, 81.1666666666667, 
    81.2083333333333, 81.25, 81.2916666666667, 81.3333333333333, 81.375, 
    81.4166666666667, 81.4583333333333, 81.5, 81.5416666666667, 
    81.5833333333333, 81.625, 81.6666666666667, 81.7083333333333, 81.75, 
    81.7916666666667, 81.8333333333333, 81.875, 81.9166666666667, 
    81.9583333333333, 82, 82.0416666666667, 82.0833333333333, 82.125, 
    82.1666666666667, 82.2083333333333, 82.25, 82.2916666666667, 
    82.3333333333333, 82.375, 82.4166666666667, 82.4583333333333, 82.5, 
    82.5416666666667, 82.5833333333333, 82.625, 82.6666666666667, 
    82.7083333333333, 82.75, 82.7916666666667, 82.8333333333333, 82.875, 
    82.9166666666667, 82.9583333333333, 83, 83.0416666666667, 
    83.0833333333333, 83.125, 83.1666666666667, 83.2083333333333, 83.25, 
    83.2916666666667, 83.3333333333333, 83.375, 83.4166666666667, 
    83.4583333333333, 83.5, 83.5416666666667, 83.5833333333333, 83.625, 
    83.6666666666667, 83.7083333333333, 83.75, 83.7916666666667, 
    83.8333333333333, 83.875, 83.9166666666667, 83.9583333333333, 84, 
    84.0416666666667, 84.0833333333333, 84.125, 84.1666666666667, 
    84.2083333333333, 84.25, 84.2916666666667, 84.3333333333333, 84.375, 
    84.4166666666667, 84.4583333333333, 84.5, 84.5416666666667, 
    84.5833333333333, 84.625, 84.6666666666667, 84.7083333333333, 84.75, 
    84.7916666666667, 84.8333333333333, 84.875, 84.9166666666667, 
    84.9583333333333, 85, 85.0416666666667, 85.0833333333333, 85.125, 
    85.1666666666667, 85.2083333333333, 85.25, 85.2916666666667, 
    85.3333333333333, 85.375, 85.4166666666667, 85.4583333333333, 85.5, 
    85.5416666666667, 85.5833333333333, 85.625, 85.6666666666667, 
    85.7083333333333, 85.75, 85.7916666666667, 85.8333333333333, 85.875, 
    85.9166666666667, 85.9583333333333, 86, 86.0416666666667, 
    86.0833333333333, 86.125, 86.1666666666667, 86.2083333333333, 86.25, 
    86.2916666666667, 86.3333333333333, 86.375, 86.4166666666667, 
    86.4583333333333, 86.5, 86.5416666666667, 86.5833333333333, 86.625, 
    86.6666666666667, 86.7083333333333, 86.75, 86.7916666666667, 
    86.8333333333333, 86.875, 86.9166666666667, 86.9583333333333, 87, 
    87.0416666666667, 87.0833333333333, 87.125, 87.1666666666667, 
    87.2083333333333, 87.25, 87.2916666666667, 87.3333333333333, 87.375, 
    87.4166666666667, 87.4583333333333, 87.5, 87.5416666666667, 
    87.5833333333333, 87.625, 87.6666666666667, 87.7083333333333, 87.75, 
    87.7916666666667, 87.8333333333333, 87.875, 87.9166666666667, 
    87.9583333333333, 88, 88.0416666666667, 88.0833333333333, 88.125, 
    88.1666666666667, 88.2083333333333, 88.25, 88.2916666666667, 
    88.3333333333333, 88.375, 88.4166666666667, 88.4583333333333, 88.5, 
    88.5416666666667, 88.5833333333333, 88.625, 88.6666666666667, 
    88.7083333333333, 88.75, 88.7916666666667, 88.8333333333333, 88.875, 
    88.9166666666667, 88.9583333333333, 89, 89.0416666666667, 
    89.0833333333333, 89.125, 89.1666666666667, 89.2083333333333, 89.25, 
    89.2916666666667, 89.3333333333333, 89.375, 89.4166666666667, 
    89.4583333333333, 89.5, 89.5416666666667, 89.5833333333333, 89.625, 
    89.6666666666667, 89.7083333333333, 89.75, 89.7916666666667, 
    89.8333333333333, 89.875, 89.9166666666667, 89.9583333333333, 90, 
    90.0416666666667, 90.0833333333333, 90.125, 90.1666666666667, 
    90.2083333333333, 90.25, 90.2916666666667, 90.3333333333333, 90.375, 
    90.4166666666667, 90.4583333333333, 90.5, 90.5416666666667, 
    90.5833333333333, 90.625, 90.6666666666667, 90.7083333333333, 90.75, 
    90.7916666666667, 90.8333333333333, 90.875, 90.9166666666667, 
    90.9583333333333, 91, 91.0416666666667, 91.0833333333333, 91.125, 
    91.1666666666667, 91.2083333333333, 91.25, 91.2916666666667, 
    91.3333333333333, 91.375, 91.4166666666667, 91.4583333333333, 91.5, 
    91.5416666666667, 91.5833333333333, 91.625, 91.6666666666667, 
    91.7083333333333, 91.75, 91.7916666666667, 91.8333333333333, 91.875, 
    91.9166666666667, 91.9583333333333, 92, 92.0416666666667, 
    92.0833333333333, 92.125, 92.1666666666667, 92.2083333333333, 92.25, 
    92.2916666666667, 92.3333333333333, 92.375, 92.4166666666667, 
    92.4583333333333, 92.5, 92.5416666666667, 92.5833333333333, 92.625, 
    92.6666666666667, 92.7083333333333, 92.75, 92.7916666666667, 
    92.8333333333333, 92.875, 92.9166666666667, 92.9583333333333, 93, 
    93.0416666666667, 93.0833333333333, 93.125, 93.1666666666667, 
    93.2083333333333, 93.25, 93.2916666666667, 93.3333333333333, 93.375, 
    93.4166666666667, 93.4583333333333, 93.5, 93.5416666666667, 
    93.5833333333333, 93.625, 93.6666666666667, 93.7083333333333, 93.75, 
    93.7916666666667, 93.8333333333333, 93.875, 93.9166666666667, 
    93.9583333333333, 94, 94.0416666666667, 94.0833333333333, 94.125, 
    94.1666666666667, 94.2083333333333, 94.25, 94.2916666666667, 
    94.3333333333333, 94.375, 94.4166666666667, 94.4583333333333, 94.5, 
    94.5416666666667, 94.5833333333333, 94.625, 94.6666666666667, 
    94.7083333333333, 94.75, 94.7916666666667, 94.8333333333333, 94.875, 
    94.9166666666667, 94.9583333333333, 95, 95.0416666666667, 
    95.0833333333333, 95.125, 95.1666666666667, 95.2083333333333, 95.25, 
    95.2916666666667, 95.3333333333333, 95.375, 95.4166666666667, 
    95.4583333333333, 95.5, 95.5416666666667, 95.5833333333333, 95.625, 
    95.6666666666667, 95.7083333333333, 95.75, 95.7916666666667, 
    95.8333333333333, 95.875, 95.9166666666667, 95.9583333333333, 96, 
    96.0416666666667, 96.0833333333333, 96.125, 96.1666666666667, 
    96.2083333333333, 96.25, 96.2916666666667, 96.3333333333333, 96.375, 
    96.4166666666667, 96.4583333333333, 96.5, 96.5416666666667, 
    96.5833333333333, 96.625, 96.6666666666667, 96.7083333333333, 96.75, 
    96.7916666666667, 96.8333333333333, 96.875, 96.9166666666667, 
    96.9583333333333, 97, 97.0416666666667, 97.0833333333333, 97.125, 
    97.1666666666667, 97.2083333333333, 97.25, 97.2916666666667, 
    97.3333333333333, 97.375, 97.4166666666667, 97.4583333333333, 97.5, 
    97.5416666666667, 97.5833333333333, 97.625, 97.6666666666667, 
    97.7083333333333, 97.75, 97.7916666666667, 97.8333333333333, 97.875, 
    97.9166666666667, 97.9583333333333, 98, 98.0416666666667, 
    98.0833333333333, 98.125, 98.1666666666667, 98.2083333333333, 98.25, 
    98.2916666666667, 98.3333333333333, 98.375, 98.4166666666667, 
    98.4583333333333, 98.5, 98.5416666666667, 98.5833333333333, 98.625, 
    98.6666666666667, 98.7083333333333, 98.75, 98.7916666666667, 
    98.8333333333333, 98.875, 98.9166666666667, 98.9583333333333, 99, 
    99.0416666666667, 99.0833333333333, 99.125, 99.1666666666667, 
    99.2083333333333, 99.25, 99.2916666666667, 99.3333333333333, 99.375, 
    99.4166666666667, 99.4583333333333, 99.5, 99.5416666666667, 
    99.5833333333333, 99.625, 99.6666666666667, 99.7083333333333, 99.75, 
    99.7916666666667, 99.8333333333333, 99.875, 99.9166666666667, 
    99.9583333333333, 100, 100.041666666667, 100.083333333333, 100.125, 
    100.166666666667, 100.208333333333, 100.25, 100.291666666667, 
    100.333333333333, 100.375, 100.416666666667, 100.458333333333, 100.5, 
    100.541666666667, 100.583333333333, 100.625, 100.666666666667, 
    100.708333333333, 100.75, 100.791666666667, 100.833333333333, 100.875, 
    100.916666666667, 100.958333333333, 101, 101.041666666667, 
    101.083333333333, 101.125, 101.166666666667, 101.208333333333, 101.25, 
    101.291666666667, 101.333333333333, 101.375, 101.416666666667, 
    101.458333333333, 101.5, 101.541666666667, 101.583333333333, 101.625, 
    101.666666666667, 101.708333333333, 101.75, 101.791666666667, 
    101.833333333333, 101.875, 101.916666666667, 101.958333333333, 102, 
    102.041666666667, 102.083333333333, 102.125, 102.166666666667, 
    102.208333333333, 102.25, 102.291666666667, 102.333333333333, 102.375, 
    102.416666666667, 102.458333333333, 102.5, 102.541666666667, 
    102.583333333333, 102.625, 102.666666666667, 102.708333333333, 102.75, 
    102.791666666667, 102.833333333333, 102.875, 102.916666666667, 
    102.958333333333, 103, 103.041666666667, 103.083333333333, 103.125, 
    103.166666666667, 103.208333333333, 103.25, 103.291666666667, 
    103.333333333333, 103.375, 103.416666666667, 103.458333333333, 103.5, 
    103.541666666667, 103.583333333333, 103.625, 103.666666666667, 
    103.708333333333, 103.75, 103.791666666667, 103.833333333333, 103.875, 
    103.916666666667, 103.958333333333, 104, 104.041666666667, 
    104.083333333333, 104.125, 104.166666666667, 104.208333333333, 104.25, 
    104.291666666667, 104.333333333333, 104.375, 104.416666666667, 
    104.458333333333, 104.5, 104.541666666667, 104.583333333333, 104.625, 
    104.666666666667, 104.708333333333, 104.75, 104.791666666667, 
    104.833333333333, 104.875, 104.916666666667, 104.958333333333, 105, 
    105.041666666667, 105.083333333333, 105.125, 105.166666666667, 
    105.208333333333, 105.25, 105.291666666667, 105.333333333333, 105.375, 
    105.416666666667, 105.458333333333, 105.5, 105.541666666667, 
    105.583333333333, 105.625, 105.666666666667, 105.708333333333, 105.75, 
    105.791666666667, 105.833333333333, 105.875, 105.916666666667, 
    105.958333333333, 106, 106.041666666667, 106.083333333333, 106.125, 
    106.166666666667, 106.208333333333, 106.25, 106.291666666667, 
    106.333333333333, 106.375, 106.416666666667, 106.458333333333, 106.5, 
    106.541666666667, 106.583333333333, 106.625, 106.666666666667, 
    106.708333333333, 106.75, 106.791666666667, 106.833333333333, 106.875, 
    106.916666666667, 106.958333333333, 107, 107.041666666667, 
    107.083333333333, 107.125, 107.166666666667, 107.208333333333, 107.25, 
    107.291666666667, 107.333333333333, 107.375, 107.416666666667, 
    107.458333333333, 107.5, 107.541666666667, 107.583333333333, 107.625, 
    107.666666666667, 107.708333333333, 107.75, 107.791666666667, 
    107.833333333333, 107.875, 107.916666666667, 107.958333333333, 108, 
    108.041666666667, 108.083333333333, 108.125, 108.166666666667, 
    108.208333333333, 108.25, 108.291666666667, 108.333333333333, 108.375, 
    108.416666666667, 108.458333333333, 108.5, 108.541666666667, 
    108.583333333333, 108.625, 108.666666666667, 108.708333333333, 108.75, 
    108.791666666667, 108.833333333333, 108.875, 108.916666666667, 
    108.958333333333, 109, 109.041666666667, 109.083333333333, 109.125, 
    109.166666666667, 109.208333333333, 109.25, 109.291666666667, 
    109.333333333333, 109.375, 109.416666666667, 109.458333333333, 109.5, 
    109.541666666667, 109.583333333333, 109.625, 109.666666666667, 
    109.708333333333, 109.75, 109.791666666667, 109.833333333333, 109.875, 
    109.916666666667, 109.958333333333, 110, 110.041666666667, 
    110.083333333333, 110.125, 110.166666666667, 110.208333333333, 110.25, 
    110.291666666667, 110.333333333333, 110.375, 110.416666666667, 
    110.458333333333, 110.5, 110.541666666667, 110.583333333333, 110.625, 
    110.666666666667, 110.708333333333, 110.75, 110.791666666667, 
    110.833333333333, 110.875, 110.916666666667, 110.958333333333, 111, 
    111.041666666667, 111.083333333333, 111.125, 111.166666666667, 
    111.208333333333, 111.25, 111.291666666667, 111.333333333333, 111.375, 
    111.416666666667, 111.458333333333, 111.5, 111.541666666667, 
    111.583333333333, 111.625, 111.666666666667, 111.708333333333, 111.75, 
    111.791666666667, 111.833333333333, 111.875, 111.916666666667, 
    111.958333333333, 112, 112.041666666667, 112.083333333333, 112.125, 
    112.166666666667, 112.208333333333, 112.25, 112.291666666667, 
    112.333333333333, 112.375, 112.416666666667, 112.458333333333, 112.5, 
    112.541666666667, 112.583333333333, 112.625, 112.666666666667, 
    112.708333333333, 112.75, 112.791666666667, 112.833333333333, 112.875, 
    112.916666666667, 112.958333333333, 113, 113.041666666667, 
    113.083333333333, 113.125, 113.166666666667, 113.208333333333, 113.25, 
    113.291666666667, 113.333333333333, 113.375, 113.416666666667, 
    113.458333333333, 113.5, 113.541666666667, 113.583333333333, 113.625, 
    113.666666666667, 113.708333333333, 113.75, 113.791666666667, 
    113.833333333333, 113.875, 113.916666666667, 113.958333333333, 114, 
    114.041666666667, 114.083333333333, 114.125, 114.166666666667, 
    114.208333333333, 114.25, 114.291666666667, 114.333333333333, 114.375, 
    114.416666666667, 114.458333333333, 114.5, 114.541666666667, 
    114.583333333333, 114.625, 114.666666666667, 114.708333333333, 114.75, 
    114.791666666667, 114.833333333333, 114.875, 114.916666666667, 
    114.958333333333, 115, 115.041666666667, 115.083333333333, 115.125, 
    115.166666666667, 115.208333333333, 115.25, 115.291666666667, 
    115.333333333333, 115.375, 115.416666666667, 115.458333333333, 115.5, 
    115.541666666667, 115.583333333333, 115.625, 115.666666666667, 
    115.708333333333, 115.75, 115.791666666667, 115.833333333333, 115.875, 
    115.916666666667, 115.958333333333, 116, 116.041666666667, 
    116.083333333333, 116.125, 116.166666666667, 116.208333333333, 116.25, 
    116.291666666667, 116.333333333333, 116.375, 116.416666666667, 
    116.458333333333, 116.5, 116.541666666667, 116.583333333333, 116.625, 
    116.666666666667, 116.708333333333, 116.75, 116.791666666667, 
    116.833333333333, 116.875, 116.916666666667, 116.958333333333, 117, 
    117.041666666667, 117.083333333333, 117.125, 117.166666666667, 
    117.208333333333, 117.25, 117.291666666667, 117.333333333333, 117.375, 
    117.416666666667, 117.458333333333, 117.5, 117.541666666667, 
    117.583333333333, 117.625, 117.666666666667, 117.708333333333, 117.75, 
    117.791666666667, 117.833333333333, 117.875, 117.916666666667, 
    117.958333333333, 118, 118.041666666667, 118.083333333333, 118.125, 
    118.166666666667, 118.208333333333, 118.25, 118.291666666667, 
    118.333333333333, 118.375, 118.416666666667, 118.458333333333, 118.5, 
    118.541666666667, 118.583333333333, 118.625, 118.666666666667, 
    118.708333333333, 118.75, 118.791666666667, 118.833333333333, 118.875, 
    118.916666666667, 118.958333333333, 119, 119.041666666667, 
    119.083333333333, 119.125, 119.166666666667, 119.208333333333, 119.25, 
    119.291666666667, 119.333333333333, 119.375, 119.416666666667, 
    119.458333333333, 119.5, 119.541666666667, 119.583333333333, 119.625, 
    119.666666666667, 119.708333333333, 119.75, 119.791666666667, 
    119.833333333333, 119.875, 119.916666666667, 119.958333333333, 120, 
    120.041666666667, 120.083333333333, 120.125, 120.166666666667, 
    120.208333333333, 120.25, 120.291666666667, 120.333333333333, 120.375, 
    120.416666666667, 120.458333333333, 120.5, 120.541666666667, 
    120.583333333333, 120.625, 120.666666666667, 120.708333333333, 120.75, 
    120.791666666667, 120.833333333333, 120.875, 120.916666666667, 
    120.958333333333, 121, 121.041666666667, 121.083333333333, 121.125, 
    121.166666666667, 121.208333333333, 121.25, 121.291666666667, 
    121.333333333333, 121.375, 121.416666666667, 121.458333333333, 121.5, 
    121.541666666667, 121.583333333333, 121.625, 121.666666666667, 
    121.708333333333, 121.75, 121.791666666667, 121.833333333333, 121.875, 
    121.916666666667, 121.958333333333, 122, 122.041666666667, 
    122.083333333333, 122.125, 122.166666666667, 122.208333333333, 122.25, 
    122.291666666667, 122.333333333333, 122.375, 122.416666666667, 
    122.458333333333, 122.5, 122.541666666667, 122.583333333333, 122.625, 
    122.666666666667, 122.708333333333, 122.75, 122.791666666667, 
    122.833333333333, 122.875, 122.916666666667, 122.958333333333, 123, 
    123.041666666667, 123.083333333333, 123.125, 123.166666666667, 
    123.208333333333, 123.25, 123.291666666667, 123.333333333333, 123.375, 
    123.416666666667, 123.458333333333, 123.5, 123.541666666667, 
    123.583333333333, 123.625, 123.666666666667, 123.708333333333, 123.75, 
    123.791666666667, 123.833333333333, 123.875, 123.916666666667, 
    123.958333333333, 124, 124.041666666667, 124.083333333333, 124.125, 
    124.166666666667, 124.208333333333, 124.25, 124.291666666667, 
    124.333333333333, 124.375, 124.416666666667, 124.458333333333, 124.5, 
    124.541666666667, 124.583333333333, 124.625, 124.666666666667, 
    124.708333333333, 124.75, 124.791666666667, 124.833333333333, 124.875, 
    124.916666666667, 124.958333333333, 125, 125.041666666667, 
    125.083333333333, 125.125, 125.166666666667, 125.208333333333, 125.25, 
    125.291666666667, 125.333333333333, 125.375, 125.416666666667, 
    125.458333333333, 125.5, 125.541666666667, 125.583333333333, 125.625, 
    125.666666666667, 125.708333333333, 125.75, 125.791666666667, 
    125.833333333333, 125.875, 125.916666666667, 125.958333333333, 126, 
    126.041666666667, 126.083333333333, 126.125, 126.166666666667, 
    126.208333333333, 126.25, 126.291666666667, 126.333333333333, 126.375, 
    126.416666666667, 126.458333333333, 126.5, 126.541666666667, 
    126.583333333333, 126.625, 126.666666666667, 126.708333333333, 126.75, 
    126.791666666667, 126.833333333333, 126.875, 126.916666666667, 
    126.958333333333, 127, 127.041666666667, 127.083333333333, 127.125, 
    127.166666666667, 127.208333333333, 127.25, 127.291666666667, 
    127.333333333333, 127.375, 127.416666666667, 127.458333333333, 127.5, 
    127.541666666667, 127.583333333333, 127.625, 127.666666666667, 
    127.708333333333, 127.75, 127.791666666667, 127.833333333333, 127.875, 
    127.916666666667, 127.958333333333, 128, 128.041666666667, 
    128.083333333333, 128.125, 128.166666666667, 128.208333333333, 128.25, 
    128.291666666667, 128.333333333333, 128.375, 128.416666666667, 
    128.458333333333, 128.5, 128.541666666667, 128.583333333333, 128.625, 
    128.666666666667, 128.708333333333, 128.75, 128.791666666667, 
    128.833333333333, 128.875, 128.916666666667, 128.958333333333, 129, 
    129.041666666667, 129.083333333333, 129.125, 129.166666666667, 
    129.208333333333, 129.25, 129.291666666667, 129.333333333333, 129.375, 
    129.416666666667, 129.458333333333, 129.5, 129.541666666667, 
    129.583333333333, 129.625, 129.666666666667, 129.708333333333, 129.75, 
    129.791666666667, 129.833333333333, 129.875, 129.916666666667, 
    129.958333333333, 130, 130.041666666667, 130.083333333333, 130.125, 
    130.166666666667, 130.208333333333, 130.25, 130.291666666667, 
    130.333333333333, 130.375, 130.416666666667, 130.458333333333, 130.5, 
    130.541666666667, 130.583333333333, 130.625, 130.666666666667, 
    130.708333333333, 130.75, 130.791666666667, 130.833333333333, 130.875, 
    130.916666666667, 130.958333333333, 131, 131.041666666667, 
    131.083333333333, 131.125, 131.166666666667, 131.208333333333, 131.25, 
    131.291666666667, 131.333333333333, 131.375, 131.416666666667, 
    131.458333333333, 131.5, 131.541666666667, 131.583333333333, 131.625, 
    131.666666666667, 131.708333333333, 131.75, 131.791666666667, 
    131.833333333333, 131.875, 131.916666666667, 131.958333333333, 132, 
    132.041666666667, 132.083333333333, 132.125, 132.166666666667, 
    132.208333333333, 132.25, 132.291666666667, 132.333333333333, 132.375, 
    132.416666666667, 132.458333333333, 132.5, 132.541666666667, 
    132.583333333333, 132.625, 132.666666666667, 132.708333333333, 132.75, 
    132.791666666667, 132.833333333333, 132.875, 132.916666666667, 
    132.958333333333, 133, 133.041666666667, 133.083333333333, 133.125, 
    133.166666666667, 133.208333333333, 133.25, 133.291666666667, 
    133.333333333333, 133.375, 133.416666666667, 133.458333333333, 133.5, 
    133.541666666667, 133.583333333333, 133.625, 133.666666666667, 
    133.708333333333, 133.75, 133.791666666667, 133.833333333333, 133.875, 
    133.916666666667, 133.958333333333, 134, 134.041666666667, 
    134.083333333333, 134.125, 134.166666666667, 134.208333333333, 134.25, 
    134.291666666667, 134.333333333333, 134.375, 134.416666666667, 
    134.458333333333, 134.5, 134.541666666667, 134.583333333333, 134.625, 
    134.666666666667, 134.708333333333, 134.75, 134.791666666667, 
    134.833333333333, 134.875, 134.916666666667, 134.958333333333, 135, 
    135.041666666667, 135.083333333333, 135.125, 135.166666666667, 
    135.208333333333, 135.25, 135.291666666667, 135.333333333333, 135.375, 
    135.416666666667, 135.458333333333, 135.5, 135.541666666667, 
    135.583333333333, 135.625, 135.666666666667, 135.708333333333, 135.75, 
    135.791666666667, 135.833333333333, 135.875, 135.916666666667, 
    135.958333333333 ;

 ycoord = 15, 25 ;

 xcoord = 10, 20, 30 ;

 Ta =
  -7.355, -7.545, -6.75, -6.6, -6.515, -6.545, -7.34, -7.17, -5.715, -3.385, 
    -2.5, -2.31, -2.12, -1.97, -1.89, -2.04, -2.135, -3.33, -4.08, -4.8, 
    -5.035, -5.04, -4.9, -5.815, -5.1, -5.15, -5.315, -5.8, -6.785, -6.35, 
    -5.995, -4.845, -0.33, 1.05, 2.065, 2.82, 3.24, 4.18, 5.065, 4.925, 
    3.445, 2.475, 0.415, -2.325, -2.92, -3.28, -3.53, -2.68, -1.465, -2.74, 
    -1.81, -1.145, -0.18, -0.495, -0.52, 0.235, 1.205, 2.535, 2.73, 3.665, 
    4.295, 4.175, 4.94, 4.9, 4.45, 4.64, 2.975, 2.725, 2.615, 2.685, 2.435, 
    1.81, 0.91, 0.205, -0.235, -0.47, -0.515, -0.64, -0.845, -1.78, -2.05, 
    -1.92, -2.125, -1.23, -1.25, -1.145, -1.6, -1.23, -1.585, -1.585, -2.3, 
    -3.15, -3.33, -3.36, -3.455, -3.855, -4.075, -4.75, -4.96, -5.165, 
    -5.515, -5.835, -6.545, -6.57, -5.72, -5.005, -4.595, -4.815, -3.385, 
    -3.49, -4.83, -4.685, -4.665, -4.815, -4.99, -5.62, -5.855, -6.195, 
    -6.57, -7.72, -6.98, -8.075, -8.33, -7.45, -7.99, -9.205, -9.06, -7.505, 
    -3.675, -0.52, -1.075, 0.005, 0.47, 0.59, 1.325, 1.63, 1.59, -0.02, 
    -1.915, -3.25, -3.25, -2.425, -4.04, -5.65, -5.835, -5.745, -5.095, 
    -5.94, -6.22, -4.83, -5.01, -4.02, 1.03, 3.93, 4.6, 4.285, 5.385, 5.39, 
    5.855, 5.045, 3.88, 2.25, -0.07, -1.25, -1.275, -1.83, -2.23, -2.965, 
    -3.6, -4.115, -3.435, -3.18, -3.76, -4.225, -3.655, -3.03, -2.51, -2.165, 
    0.25, 0.005, 0.1, -0.37, -0.09, 0.575, -0.515, -1.49, -1.795, -1.965, 
    -2.835, -2.945, -2.88, -3.1, -3.305, -3.18, -3.02, -3.015, -2.87, -2.635, 
    -2.615, -2.5, -2.25, -1.475, -1.045, -0.975, -0.885, -0.44, 0.04, 0.575, 
    0.585, 0.22, -0.6, -1.41, -1.905, -2.355, -2.885, -3.295, -3.56, -3.7, 
    -3.8, -4.255, -4.765, -5.17, -5.03, -5.185, -4.64, -3.875, -3.515, 
    -1.445, -0.825, -1.09, -1.695, -2.995, -3.1, -3.2, -3.325, -3.35, -3.39, 
    -3.75, -3.445, -3.285, -3.715, -4.055, -3.645, -3.545, -3.24, -2.81, 
    -2.575, -2.42, -2.11, -1.765, -1.535, -1.51, -1.54, -1.775, -1.7, -0.625, 
    -0.39, -0.87, -1.65, -2.055, -2.42, -2.41, -2.55, -2.84, -2.545, -2.04, 
    -2.205, -2.17, -2.405, -3.215, -3.525, -3.61, 0.655, 3.6, 5.785, 6.57, 
    6.995, 7.15, 7.53, 7.385, 5.8, 4.335, 4.11, 4.4, 4.24, 4.335, 4.73, 
    4.535, 2.89, 1.555, 0.325, 0.35, 0.845, 0.995, 0.935, 1.355, 1.905, 
    4.155, 4.245, 4.125, 6.345, 5.6, 5.915, 5.98, 5.43, 4.75, 4.135, 3.435, 
    1.83, 1.76, 2.32, 1.64, 0.425, 0.01, -0.145, -0.32, -0.23, -0.18, -0.03, 
    0.285, 0.6, 1.02, 1.555, 2.43, 3, 4.035, 3.705, 3.68, 3.845, 3.64, 2.905, 
    3.01, 3.07, 3.265, 3.21, 2.86, 2.855, 2.865, 2.67, 2.83, 2.345, 1.865, 
    1.64, 1.73, 3.605, 3.61, 3.465, 3.61, 4.065, 4.53, 5.265, 5.195, 5.21, 
    4.105, 3.33, 3.12, 2.525, 1.895, 0.15, 1.09, 0, -0.015, -0.63, 0.365, 
    0.835, -0.315, -0.39, -0.23, 4.315, 6.37, 6.895, 7.54, 8.86, 9.645, 
    9.965, 10.18, 9.68, 7.155, 4.065, 3.22, 3.015, 2.745, 2.37, 2.38, 2.035, 
    2.295, 1.67, 3.37, 4.295, 3.935, 3.145, 3.32, 8.21, 11.115, 11.675, 
    12.655, 13.19, 13.435, 13.86, 13.49, 12.665, 10.17, 7.065, 5.96, 5.635, 
    5.365, 5.86, 5.51, 6.28, 7.3, 6.65, 6.65, 6.48, 6.695, 5.76, 5.82, 10.15, 
    11.875, 13.14, 14.395, 14.8, 14.755, 14.34, 14.805, 13.355, 10.935, 
    8.645, 7.925, 8.335, 8.8, 9.5, 9.395, 9.405, 9.295, 9.275, 8.95, 8.11, 
    6.99, 5.58, 2.68, 3.73, 6.09, 8.08, 7.55, 8.205, 8.445, 7.735, 7.105, 
    3.555, 1.365, 1.605, 0.555, -0.095, -0.245, -0.26, -0.435, -0.365, 
    -0.355, -0.08, -0.255, -0.205, -0.09, -0.065, -0.125, -0.135, 0.01, 
    1.385, 1.325, 2.04, 1.44, 0.56, 1.59, 2, 0.745, -0.065, -1.02, -1.85, 
    -2.13, -2.685, -2.695, -2.875, -2.955, -3.25, -3.665, -3.755, -3.6, 
    -3.76, -3.7, -0.905, -0.065, 1.235, 1.45, 1.37, 1.02, 2.045, 3.05, 2.44, 
    0.715, 0.185, -0.005, -0.605, -0.89, -0.365, -0.47, -0.855, -0.65, 
    -0.475, -0.29, -0.12, -0.145, -1.565, -1.24, -0.695, 0.885, 3.405, 3.905, 
    4.145, 5.08, 5.135, 4.29, 3.015, 1.875, 1.085, 0.55, 0.14, -0.35, -0.775, 
    -1.04, -1.3, -1.82, -2.17, -1.585, -2.265, -1.475, -1.1, -0.55, -0.065, 
    0.42, 1.105, 1.775, 1.865, 1.84, 1.32, 1.39, 1.325, 1.255, 0.875, 1.505, 
    1.655, 0.38, -0.1, -0.275, -0.385, -0.22, 0.45, 0.43, 0.49, 0.57, 0.58, 
    0.53, 0.44, 0.31, 0.385, 0.665, 1.135, 0.99, 1.275, 0.67, 0.04, -1.21, 
    -2.36, -3.435, -3.77, -4.13, -4.62, -4.36, -5.16, -5.175, -5.795, -6.895, 
    -7.15, -7.68, -8.83, -8.525, -5.37, -3.675, -2.575, -2.4, -1.495, -1.24, 
    -1.025, -0.9, -1.645, -3.29, -4.665, -5.31, -6.23, -6.83, -6.85, -6.555, 
    -6.935, -6.27, -5.78, -4.76, -4.385, -5.055, -4.825, -4.195, -2.995, 
    -0.53, 0.425, 0.46, 1.77, 2.12, 1.37, 1.625, 0.675, -0.295, -0.265, 0.47, 
    0.575, 0.845, 1.185, 2.2, 1.26, -1.705, -3.45, -4.61, -5.7, -7.2, -7.61, 
    -7.88, -8.115, -8.325, -8.22, -6.61, -5.275, -5.45, -5.67, -7.43, -8.115, 
    -9.05, -9.905, -9.425, -9.425, -9.975, -10.41, -10.37, -10.525, -10.585, 
    -10.59, -10.185, -10.37, -10.9, -10.375, -10.3, -9.47, -7.345, -4.955, 
    -4.905, -4.81, -3.835, -3.385, -4.11, -4.87, -6.115, -6.84, -7.425, 
    -7.925, -8.435, -8.58, -8.355, -8.895, -9.32, -10.21, -11.555, -10.74, 
    -9.74, -11.12, -11.795, -8.96, -8.105, -6.325, -5.97, -5.05, -4.475, 
    -5.55, -6.345, -7.165, -8.095, -8.82, -9.12, -9.48, -9.46, -9.425, 
    -9.385, -9.26, -8.82, -8.485, -8.135, -7.27, -6.12, -5.78, -4.615, 
    -3.995, -4.02, -4.47, -3.84, -3.655, -3.445, -2.9, -2.355, -2.185, 
    -2.095, -1.985, -1.8, -1.595, -1.53, -1.515, -1.49, -1.565, -1.435, 
    -1.435, -1.68, -1.955, -2.365, -2.435, -2.37, -1.365, -0.055, 0.575, 1.5, 
    3.035, 3.68, 4.335, 4.95, 3.63, 1.775, 0.865, 0.36, 0.275, 0.995, 1.82, 
    1.785, 1.4, 1.36, 1.285, 1.6, 1.835, 1.875, 1.515, 1.73, 3.245, 4.875, 
    5.565, 6.04, 5.82, 5.32, 5.02, 4.055, 4.01, 3.235, 2.145, 1.935, 1.62, 
    1.66, 1.345, 1.35, 0.745, 0.8, 0.725, 0.695, 0.09, 0.1, -0.44, -0.665, 
    1.735, 4.885, 5.61, 6.485, 6.69, 6.055, 6.27, 5.845, 5.125, 3.245, 1.01, 
    0.41, 1.095, 0.325, 0.5, 0.305, 0.655, 1.325, 1.02, 1.255, 0.355, 0.56, 
    0.72, 0.96, 3.15, 5.19, 5.59, 7.01, 7.335, 7.925, 7.875, 7.895, 6.835, 
    4.98, 2.54, 0.655, 0.6, 0.4, 0.27, 0.49, 0.76, 0.82, 1.415, 3.575, 4.175, 
    1.61, 1.81, 1.805, 5.895, 10.93, 11.875, 12.64, 13.65, 14.125, 14.33, 
    13.455, 11.69, 8.375, 6.52, 6.475, 8.25, 8.96, 7.66, 7.7, 7.52, 7.625, 
    7.815, 6.98, 4.965, 3.055, 2.155, 4.905, 7.49, 9.84, 11.135, 12.03, 
    12.36, 11.785, 12.515, 10.92, 10.01, 8.255, 7.295, 6.835, 7.165, 7.89, 
    8.21, 7.47, 6.67, 6.075, 6.055, 5.65, 5.05, 4.79, 4.53, 4.405, 4.635, 
    6.24, 6.61, 6.805, 7.015, 6.83, 6.02, 4.875, 4.105, 3.2, 2.305, 2.36, 
    2.155, 1.6, 1.145, 0.875, 0.415, -0.01, -0.35, -0.21, -0.37, -0.445, 
    -0.4, -0.04, 0.475, 2.315, 3.425, 4.885, 5.01, 3.305, 2.65, 1.91, 2.11, 
    1.01, -0.785, -2.23, -2.46, -2.97, -3.2, -2.71, -2.51, -2.93, -3.775, 
    -4.095, -4.535, -4.84, -6.07, -6.715, -3.515, -0.39, -0.05, -0.225, 0.32, 
    0.97, 1.155, 0.89, 0.04, -2.045, -3.91, -4.535, -4.6, -5.05, -5.16, 
    -4.72, -4.505, -5.255, -6.435, -6.42, -5.605, -5.01, -5.03, -4.77, 
    -2.195, 2.48, 4.08, 5.16, 5.565, 5.865, 6.11, 5.7, 4.06, 1.125, 0.435, 
    1.28, 0.965, 0.3, 1.215, 0.53, 0.51, 1.36, 0.055, -0.23, -0.62, 0, 0.895, 
    0.905, 1.045, 2.225, 3.185, 4.6, 4.88, 5.415, 4.655, 4.425, 3.8, 1.905, 
    -0.445, -1.38, -1.93, -1.92, 0.985, 2.22, 2.435, 1.735, 1.81, 2.32, 
    2.415, 1.915, 0.91, 2.285, 2.85, 5.575, 7.23, 8.69, 8.46, 7.6, 6.61, 6.31, 
    6.02, 5.235, 4.925, 4.94, 4.37, 3.765, 5.105, 5.15, 4.895, 4.455, 3.955, 
    3.905, 3.905, 3.665, 3.23, 2.34, 2.375, 2.05, 0.97, 0.635, -1.855, -2.95, 
    -3.085, -3.63, -4.23, -5.015, -5.825, -6.425, -7.33, -8.405, -8.91, 
    -8.615, -9.645, -10.04, -10.88, -11.45, -11.965, -12.235, -12.515, 
    -12.415, -10.93, -8.25, -6.695, -6.955, -5.96, -7.365, -6.795, -7.075, 
    -7.945, -9.305, -11.035, -11.44, -11.825, -11.58, -12.035, -12.755, 
    -12.61, -11.075, -10.5, -10.245, -9.655, -9.535, -9.825, -9.65, -9.095, 
    -8.31, -7.095, -7.035, -6.855, -7.495, -8.515, -9.36, -9.965, -10.825, 
    -11.33, -11.56, -11.925, -12.32, -12.825, -12.88, -13.815, -14.32, 
    -14.955, -14.53, -14.415, -14.87, -14.375, -14.77, -14.145, -10.085, 
    -9.09, -8.33, -6.735, -7.955, -7.56, -8.015, -9.275, -10.56, -12.09, 
    -12.675, -13.005, -12.425, -11.535, -10.825, -10.895, -10.755, -10.785, 
    -10.695, -10.23, -10.43, -10.04, -9.725, -7.485, -1.285, -0.29, -0.16, 
    -0.38, -0.045, -0.255, 0.37, -1.49, -2.965, -3.435, -3.87, -3.155, 
    -2.305, -2.33, -2.59, -2.8, -1.925, -1.735, -1.4, -2.195, -2.29, -0.96, 
    -2.005, 0.03, 5.11, 6.15, 6.175, 7.57, 7.14, 7.885, 6.83, 4.14, 0.645, 
    -0.96, -0.375, -0.04, -0.23, -0.145, -0.28, -1.02, 0.615, 0.77, 0.62, 
    0.16, 0.315, -0.91, -2.27, -0.615, 4.14, 4.54, 3.83, 3.195, 3.43, 3.36, 
    2.745, 0.845, -0.315, -1.91, -2.33, -2.745, -3.535, -4.07, -5.01, -5.47, 
    -5.905, -7.04, -7.385, -7.685, -7.2, -6.375, -6.535, -5.69, -3.28, 
    -0.525, 0.79, 0.905, 1.02, 1.56, 1.49, -0.495, -2.175, -2.895, -3.095, 
    -3.4, -2.645, -1.965, -2.055, -2.165, -2.97, -4.335, -3.815, -2.18, 0.21, 
    0.665, 0.43, 0.655, 3.58, 3.495, 4.245, 4.465, 4.85, 4.59, 4.26, 3.67, 
    2.045, 1.785, 2.055, 2.625, 2.445, 2.395, 2.105, 1.475, 0.92, -0.795, 
    -2.14, -3.39, -5.35, -5.66, -5.84, -6.37, -6.355, -6.04, -6.16, -6.745, 
    -6.245, -6.955, -7.37, -8, -8.72, -9.125, -9.62, -10.505, -11.24, -11.81, 
    -12.43, -12.6, -13.06, -13.38, -11.865, -10.825, -10.53, -11.27, -10.905, 
    -9.55, -7.595, -4.085, -3.155, -4.43, -5.375, -6.38, -6.51, -6.2, -7.65, 
    -8.285, -8.77, -9.165, -9.735, -10.02, -10.195, -10.51, -10.71, -10.93, 
    -11.065, -11, -11.06, -11.17, -11.32, -11.375, -10.61, -9.92, -8.895, 
    -8.965, -8.75, -8.755, -9.17, -10.595, -10.675, -10.62, -11.175, -11.345, 
    -11.39, -11.695, -11.66, -11.335, -11.495, -12.24, -12.115, -12.18, 
    -12.14, -11.995, -11.935, -10.885, -7.475, -4.39, -2.31, -2.73, -2.565, 
    -1.045, -1.31, -3.53, -4.64, -4.62, -4.335, -5.515, -5.86, -5.425, 
    -5.865, -5.865, -5.38, -5.42, -5.465, -5.11, -4.655, -5, -5.305, -3.68, 
    0.3, 1.87, 2.7, 3.505, 3.69, 4.08, 3.49, 1.735, -0.97, -2.08, -2.675, 
    -3.06, -3.27, -3.89, -3.07, -1.875, -2.305, -2.15, -2.1, -2.715, -2.985, 
    -0.955, -0.215, 0.515, 5.195, 8.785, 9.225, 8.35, 8.725, 7.705, 6.05, 
    3.71, 0.975, -1.16, -2.095, -1.58, -1.835, -0.91, -0.03, -1.605, -1.17, 
    -1.895, -1.175, -1.545, -2.025, -3.73, -3.86, -3.345, 2.315, 3.785, 
    5.015, 4.19, 3.585, 3.145, 2.52, 1.955, -1.575, -3.39, -3.575, -3.205, 
    -2.665, -2.745, -2.525, -2.835, -2.58, -2.665, -2.57, -3.01, -3.335, 
    -3.565, -3.855, -3.535, -2.955, -1.765, 0.75, 1.5, 1.08, 0.455, 0.315, 
    -1.165, -2.665, -3.43, -4.005, -4.715, -5.455, -5.78, -6.79, -7.465, 
    -7.335, -7.735, -7.89, -6.925, -6.36, -5.835, -6.605, -6.105, -2.23, 
    -0.71, 0.665, 1.175, 1.4, 1.33, 0.61, -1.795, -3.185, -4.505, -5.175, 
    -5.71, -6.015, -5.5, -5.5, -5.585, -5.24, -4.56, -4.76, -4.69, -4.35, 
    -4.465, -4.26, -3.565, 1.83, 3.505, 2.76, 2.385, 2.26, 2.495, 1.51, 
    0.325, -1.195, -1.64, -2.145, -2.565, -3.025, -3.54, -3.24, -3.705, 
    -4.01, -4.6, -4.815, -4.81, -4.86, -5.15, -5.755, -5.32, -3.705, -2.425, 
    -1.77, -2.05, -3.41, -4.075, -4.72, -5.075, -5.605, -6.04, -6.7, -7.5, 
    -7.795, -8.12, -8.675, -10.235, -11.22, -11.485, -12.015, -12.63, -13.78, 
    -15.085, -15.58, -14.845, -11.125, -8.695, -6.685, -6.2, -6.495, -6.385, 
    -7.42, -9.66, -11.865, -13.28, -14.14, -14.65, -15.61, -16.54, -16.78, 
    -17.69, -17.96, -18.28, -18.675, -19.345, -19.56, -19.125, -19.805, 
    -19.305, -14.49, -11.81, -11.34, -11.38, -10.775, -10.575, -10.95, 
    -12.405, -14.26, -15.32, -16.83, -15.885, -16.525, -16.755, -16.51, 
    -15.7, -15.335, -15.35, -15.14, -14.785, -14.17, -13.585, -13.835, 
    -14.24, -12.725, -10.805, -9.535, -7.9, -7.18, -6.33, -7.795, -9.215, 
    -10.115, -9.975, -9.47, -9.36, -9.225, -8.995, -9.485, -9.485, -9.63, 
    -10.185, -11.245, -9.905, -9.77, -10.84, -12.165, -12.645, -12.71, 
    -12.485, -11.98, -10.905, -10.755, -11.565, -12.84, -14.165, -15.435, 
    -15.755, -15.655, -16.355, -17.17, -16.77, -16.02, -15.865, -16.38, 
    -17.825, -18.595, -19.02, -19.315, -19.555, -19.755, -19.985, -19.705, 
    -19.19, -18.81, -18.725, -18.26, -18.495, -18.97, -19.66, -20.705, 
    -21.335, -21.745, -22.295, -23.25, -24.245, -24.665, -24.505, -24.485, 
    -24.37, -24.205, -23.345, -22.25, -22.24, -22.17, -22.07, -21.72, 
    -18.895, -19.35, -17.555, -14.885, -12.675, -15.025, -18.625, -17.785, 
    -16.245, -17.095, -16.09, -16.875, -17.51, -18.045, -18.28, -18.3, 
    -18.415, -17.535, -16.975, -17.025, -17.1, -17.755, -18.285, -18.105, 
    -18.125, -17.525, -17.12, -17.48, -18.1, -18.54, -19.775, -20.585, 
    -21.17, -21.385, -21.095, -21.08, -21.235, -20.99, -20.805, -20.515, 
    -20.42, -20.185, -20.075, -20.405, -20.71, -21.015, -20.97, -20.575, 
    -20.225, -19.76, -19.475, -19.22, -19.465, -19.27, -19.115, -19.405, 
    -19.44, -19.37, -19.37, -19.395, -19.415, -19.415, -19.275, -19.17, 
    -19.21, -19.08, -18.99, -18.95, -18.815, -19.28, -18.905, -15.135, 
    -12.275, -11.595, -10.325, -10.455, -11.855, -12.435, -14.485, -15.87, 
    -17.055, -16.975, -16.375, -16.115, -16.07, -16, -15.48, -15.11, -14.535, 
    -14.875, -14.745, -14.215, -13.755, -13.425, -12.825, -10.51, -7.39, 
    -5.575, -4.445, -4.69, -4.975, -6.65, -7.895, -9.725, -11.065, -10.655, 
    -11.37, -10.1, -9.975, -9.885, -9.42, -9.41, -8.945, -8.61, -8.47, 
    -8.175, -7.835, -7.43, -7.385, -7.315, -6.92, -6.52, -6.23, -5.77, -5.79, 
    -6.225, -6.285, -6.125, -5.98, -5.755, -5.645, -5.51, -5.42, -5.425, 
    -5.535, -5.615, -5.5, -5.315, -5.195, -5.08, -5.12, -5.225, -5.365, 
    -5.59, -5.365, -5.44, -5.41, -5.505, -5.91, -6.135, -6.27, -6.38, -6.515, 
    -6.58, -6.55, -6.56, -6.645, -6.965, -7.265, -7.38, -7.825, -7.89, -7.78, 
    -7.7, -7.755, -7.95, -8.075, -8.12, -8.325, -8.255, -7.81, -8.43, -8.73, 
    -8.65, -9.255, -9.505, -9.465, -9.515, -9.92, -10.06, -10.07, -10.025, 
    -9.935, -9.81, -9.62, -8.785, -8.325, -8.485, -8.735, -8.785, -8.92, 
    -5.815, -4.445, -2.155, -2.13, -4.205, -4.08, -5.545, -6.225, -6.72, 
    -6.51, -6.09, -5.84, -5.775, -5.79, -5.185, -5.145, -4.935, -4.48, -4.06, 
    -3.765, -3.84, -4.545, -4.635, -3.765, -2.795, -2.095, -2.21, -2.855, 
    -3.545, -3.3, -3.06, -2.925, -3.525, -3.695, -3.95, -3.685, -3.495, 
    -3.18, -2.925, -3.41, -3.555, -3.325, -3.215, -3.42, -3.67, -3.945, 
    -4.09, -4.305, -4.125, -3.16, -3.65, -3.36, -2.73, -2.61, -3.21, -4.645, 
    -5.35, -5.675, -5.55, -5.51, -5.575, -5.635, -6.055, -6.94, -7.69, 
    -8.405, -9.185, -8.205, -7.705, -7.895, -7.725, -7.58, -6.49, -3.005, 
    -4.335, -3.93, -4.2, -3.965, -5.115, -6.095, -7.21, -7.88, -8.145, 
    -8.285, -8.885, -8.875, -8.96, -9.115, -8.93, -9.305, -9.47, -9.33, 
    -7.835, -7.315, -7.565, -7.18, -6.55, -5.3, -4.76, -4.48, -4.66, -4.61, 
    -4.58, -4.835, -5.255, -5.445, -5.325, -5.35, -5.245, -5.005, -4.79, 
    -4.74, -4.655, -4.06, -3.845, -3.125, -3.29, -2.995, -3.185, -3.31, 
    -2.025, 1.175, 2.505, 3.175, 3.145, 2.57, 1.095, -1.35, -2.875, -3.63, 
    -4.415, -5.305, -5.74, -4.94, -4.63, -4.425, -4.875, -5.035, -4.79, 
    -5.865, -5.805, -5.955, -5.34, -5.38, -2.91, -0.385, -0.27, 0.215, -0.42, 
    -0.215, -1.255, -2.87, -4.465, -5.465, -7.125, -7.495, -6.945, -5.57, 
    -5.24, -4.35, -4.25, -4.575, -4.62, -4.525, -4.58, -5.09, -5.075, -5.31, 
    -5.065, -4.22, -4.815, -5.265, -5.525, -6.25, -6.02, -6.115, -6.55, 
    -6.92, -6.215, -5.89, -5.82, -5.755, -5.795, -6.735, -8.43, -9.43, -8.76, 
    -8.13, -7.59, -7.745, -8.195, -8.035, -7.89, -7.93, -8.515, -8.45, -8.89, 
    -9.35, -10.29, -11.62, -12.92, -13.94, -14.675, -15.21, -16, -16.61, 
    -16.38, -17.19, -17.32, -17.855, -17.57, -18.915, -18.505, -17.815, 
    -18.93, -19.07, -15.53, -13.015, -12.67, -12.56, -12.655, -11.455, 
    -12.965, -14.29, -15.45, -15.815, -15.785, -15.355, -14.63, -14.145, 
    -14.09, -14.285, -14.1, -13.745, -13.875, -14.36, -14.435, -13.25, -12.4, 
    -12.58, -11.29, -8.965, -8.625, -8.975, -9.55, -10.125, -11.08, -11.315, 
    -12.695, -13.315, -13.875, -13.795, -14.37, -14.84, -13.87, -13.465, 
    -13.915, -14.755, -15.205, -15.305, -15.57, -15.355, -15.43, -14.65, 
    -9.12, -4.545, -3, -5.655, -6.365, -6.82, -6.97, -8.125, -10.44, -12.505, 
    -12.785, -12.57, -11.98, -11.945, -12.24, -11.8, -11.285, -10.035, 
    -10.09, -9.615, -10.11, -10.335, -9.92, -10.165, -7.91, -5.725, -5.41, 
    -5.31, -5.18, -5.97, -6.53, -7.595, -8.935, -9.815, -10.375, -10.545, 
    -11.495, -11.895, -12.705, -12.995, -12.85, -13.365, -12.865, -13.145, 
    -13.335, -13.625, -11.99, -12.155, -7.805, -2.85, -2.62, -2.51, -2.495, 
    -2.89, -3.86, -5.75, -8.58, -10.49, -9.89, -9.2, -9.57, -9.025, -9.41, 
    -9.21, -10.37, -10.85, -10.56, -9.405, -9.39, -10.125, -10.545, -9.535, 
    -8.555, -7.765, -8.935, -8.975, -8.225, -8.225, -8.305, -9.36, -10.3, 
    -10.46, -10.32, -10.325, -10.44, -10.57, -10.73, -10.81, -10.83, -10.85, 
    -10.68, -10.515, -10.485, -10.46, -10.375, -10.2, -9.87, -9.71, -9.97, 
    -10.115, -10.29, -10.265, -10.525, -10.655, -10.83, -11.13, -11.32, 
    -11.45, -11.365, -11.41, -11.175, -11, -11.05, -11.16, -11.21, -11.25, 
    -11.325, -11.46, -11.74, -11.78, -11.23, -10.245, -9.775, -9.115, -8.925, 
    -10.265, -10.64, -11.025, -11.22, -11.205, -11.165, -11, -10.64, -10.21, 
    -9.67, -8.725, -7.44, -7.26, -7.165, -6.45, -6.07, -5.98, -5.965, -5.635, 
    -4.63, -3.835, -3.85, -3.82, -4.06, -3.585, -4.02, -4.765, -5.095, -5.26, 
    -5.36, -5, -4.545, -4.355, -4.075, -4.35, -4.48, -4.435, -4.39, -4.57, 
    -4.73, -5.175, -5.51, -6.235, -6.595, -6.35, -6.12, -6.375, -5.735, 
    -6.26, -6.19, -6.82, -7.175, -7.385, -7.775, -8.295, -8.16, -8.425, 
    -8.16, -7.82, -7.76, -7.835, -7.975, -8.065, -8.135, -8.09, -7.875, 
    -7.91, -7.56, -6.925, -5.675, -5.265, -4.71, -4.275, -5.165, -7.075, 
    -7.53, -8.385, -10.07, -11.04, -9.97, -9.465, -9.525, -9.72, -9.175, 
    -8.805, -9.18, -8.68, -9.065, -9.46, -9.745, -8.465, -6.73, -3.945, 
    -0.485, -0.495, -0.645, -2.17, -4.61, -5.76, -6.04, -6.25, -6.28, -5.96, 
    -6.185, -5.615, -5.485, -5.62, -5.33, -5.25, -5.07, -4.695, -4.665, 
    -4.62, -4.345, -4.385, -4.2, -4.09, -4.535, -3.27, -3.08, -3.26, -3.99, 
    -4.615, -5.075, -5.045, -4.375, -4.35, -4.355, -4.49, -4.785, -4.645, 
    -4.725, -4.53, -4.265, -4.075, -3.99, -3.95, -3.695, -3.64, -3.775, 
    -3.84, -3.81, -3.76, -3.865, -4.39, -4.74, -5.52, -6.44, -7.42, -7.99, 
    -8.725, -10.68, -12.035, -12.77, -12.49, -13.635, -15.155, -15.77, 
    -16.06, -16.15, -15.66, -15.92, -15.74, -12.88, -9.905, -6.055, -4.78, 
    -5.285, -5.765, -7.07, -8.32, -10.375, -12.445, -12.86, -12.95, -13.015, 
    -12.6, -12.31, -11.595, -11.38, -11.495, -11.11, -11.01, -10.505, -10.46, 
    -10.64, -10.375, -7.355, -3.06, -0.025, 0.585, -1.085, -1.615, -2.14, 
    -2.935, -4.09, -4.345, -5.01, -4.615, -4.715, -4.73, -4.525, -4.585, 
    -4.71, -5.085, -4.83, -4.06, -4.135, -4.375, -4.645, -5.415, -4.645, 
    -2.545, -1.125, -0.895, -0.94, -1.635, -2.395, -2.705, -3.54, -4.98, 
    -4.475, -4.38, -4.09, -5.535, -5.845, -5.85, -4.81, -4.02, -4.13, -4.63, 
    -5.645, -5.195, -5.64, -5.865, -2.765, 0.66, 1.53, 1.22, 1.9, 1.68, 1.07, 
    -0.37, -1.655, -3.4, -4.36, -4.665, -4.765, -4.8, -4.94, -5.55, -5.315, 
    -5.13, -4.915, -5.165, -5.695, -5.65, -5.645, -5.63, -1.34, 2.43, 3.78, 
    4.19, 3.38, 3.8, 3.395, 1.47, 0.345, -0.085, -0.675, -0.12, -2.305, 
    -4.25, -4.78, -4.225, -4.34, -5.215, -5.575, -2.12, -3.445, -1.35, 
    -0.435, -0.095, 1.43, 1.76, 2.09, 2.54, 2.19, 1.905, 1.185, 1.175, 
    -0.655, -1.435, -2.045, -1.88, -3.135, -3.9, -3.785, -2.76, -2.755, 
    -2.575, -3.11, -4.3, -5.945, -6.455, -6.14, -5.77, -3.155, 0.405, 2.715, 
    2.23, 2.61, 0.42, 1.26, -0.115, -1.685, -2.155, -2.805, -3.24, -3.125, 
    -3.45, -4.3, -4.965, -5.03, -5.665, -5.7, -5.585, -5.795, -5.925, -6.055, 
    -6.155, -5.78, -5.09, -5.12, -4.5, -4.32, -4.195, -4.57, -5.32, -6.03, 
    -6.63, -7.41, -8.055, -8.335, -8.65, -8.58, -8.6, -9.29, -10.37, -10.12, 
    -9.49, -8.435, -8.325, -9.545, -7.535, -6.17, -4.84, -3.28, -2.545, 
    -2.07, -1.18, -1.835, -2.55, -2.56, -2.47, -2.72, -2.68, -3.175, -3.03, 
    -2.35, -2.535, -3.365, -3.07, -3.2, -3.105, -4.345, -3.715, -3.79, 
    -3.585, -1.015, 0.52, 2.87, 3.41, 2.845, 1.565, 1.67, 0.03, -2.025, 
    -2.87, -3.785, -3.61, -3.735, -3.275, -2.905, -3.425, -2.73, -3.705, 
    -3.81, -4.375, -5.085, -6.665, -5.465, -4.25, -1.75, 1.065, 0.805, 1.4, 
    2.235, 2.115, 1.685, -0.19, -2.595, -4.095, -4.015, -3.665, -3.205, 
    -3.03, -2.985, -3.485, -4.155, -4.565, -5.53, -5.695, -4.95, -5.59, 
    -5.92, -5.84, -5.445, -4.705, -4.615, -3.24, -3.86, -3.725, -4.13, -4.04, 
    -4.295, -4.435, -4.19, -4.33, -4.815, -5.005, -5.065, -4.825, -4.8, 
    -4.64, -4.24, -4.485, -4.825, -4.995, -5.245, -5.265, -5.22, -5.775, 
    -5.79, -5.325, -4.55, -5.65, -5.77, -5.91, -7.145, -7.855, -9.365, -8.31, 
    -7.795, -7.275, -7.145, -7.52, -7.775, -7.36, -7.85, -8.25, -8.15, -8.14, 
    -8.6, -8.595, -7.36, -5.85, -4.705, -5.065, -5.045, -5.975, -5.795, 
    -5.55, -6.68, -7.605, -8.11, -7.86, -7.685, -7.485, -7.135, -7.315, 
    -7.36, -7.205, -6.965, -6.82, -6.835, -6.99, -6.895, -6.84, -6.525, 
    -6.02, -5.675, -4.24, -4.675, -4.665, -4.695, -5.27, -6.405, -7.235, 
    -7.1, -7.345, -7.725, -7.48, -7.275, -7.79, -7.68, -7.6, -7.385, -6.56, 
    -5.955, -6.11, -6.545, -6.635, -6.515, -6.17, -5.305, -5.655, -6.005, 
    -6.695, -7.035, -7.16, -7.205, -7.37, -7.59, -7.7, -7.82, -8.26, -8.495, 
    -8.565, -8.605, -8.81, -9.19, -9.41, -9.475, -9.51, -9.555, -9.64, -9.5, 
    -9.35, -9.2, -9.22, -9.44, -9.615, -9.78, -9.78, -9.685, -9.65, -9.625, 
    -9.6, -9.625, -9.74, -9.875, -9.965, -10.075, -10.175, -10.23, -10.215, 
    -10.255, -10.31, -10.31, -10.375, -10.22, -9.755, -8.63, -7.215, -8.505, 
    -9.28, -9.46, -10.105, -10.5, -10.91, -11.29, -11.585, -11.655, -11.925, 
    -12.14, -12.165, -11.54, -11.055, -11.17, -11.26, -10.815, -10.49, 
    -10.505, -10.025, -9.39, -9.115, -8.83, -8.345, -6.725, -6.045, -5.165, 
    -5.88, -7.2, -7.63, -7.795, -8.485, -10.6, -11.19, -9.17, -8.75, -9.605, 
    -10.255, -10.735, -10.06, -8.325, -6.455, -6.355, -6.43, -5.34, -3.955, 
    -2.875, -3.755, -3.085, -2.67, -2.3, -3.165, -4.445, -5.105, -5.345, 
    -5.525, -6.06, -6.5, -7.16, -7.35, -7.11, -8.16, -8.68, -8.495, -8.6, 
    -8.165, -7.945, -8.435, -6.715, -4.175, -2.98, -2.245, -2.635, -2.99, 
    -3.59, -4.015, -5.26, -6.64, -6.955, -6.945, -6.925, -6.8, -7.245, -7.65, 
    -8, -8.105, -8.07, -7.99, -8.055, -8.935, -9.44, -9.425, -6.345, -4.485, 
    -3.795, -3.12, -2.88, -2.25, -2.125, -3.3, -5.79, -7.66, -8.255, -8.985, 
    -9.48, -9.625, -10.43, -10.325, -9.5, -10.63, -10.7, -10.325, -10.52, 
    -10.815, -10.675, -10.165, -6.18, -3.14, -1.37, -1.145, -0.9, -0.62, 
    -0.66, -3.105, -4.88, -6.73, -6.945, -7.765, -8.805, -8.975, -8.825, 
    -8.2, -7.88, -9.39, -8.385, -8.9, -7.305, -7.37, -9.75, -9.985, -6.56, 
    -1.025, 1.22, 1.44, 0.785, 0.615, 0.5, -1.65, -3.605, -4.805, -5.71, 
    -5.435, -5.24, -5.53, -5.61, -5.725, -6.06, -6.46, -6.985, -7.275, 
    -7.265, -7.285, -7.25, -7.255, -7.085, -6.685, -6.695, -6.635, -6.77, 
    -6.92, -6.815, -7.225, -7.32, -7.365, -7.32, -7.345, -7.475, -7.72, 
    -7.725, -7.9, -8.01, -8.005, -8.005, -8.155, -8.295, -8.405, -8.615, 
    -8.675, -8.375, -7.33, -6.57, -6.145, -7.515, -6.66, -5.42, -6.335, 
    -7.645, -8.825, -9.915, -11.955, -11.91, -11.31, -10.255, -10.925, 
    -10.965, -10.295, -9.375, -9.245, -9.375, -9.755, -10.95, -10.68, -6.425, 
    -0.755, -0.125, -1.15, -2.785, -3.34, -3.385, -3.89, -4.725, -6.705, 
    -7.995, -7.465, -7.3, -7.64, -9.24, -9.84, -10.31, -9.99, -9.83, -9.6, 
    -9.3, -8.495, -7.625, -6.185, -4.885, -5.4, -4.21, -1.24, -1.065, -1.255, 
    -1.425, -2.215, -3.815, -5.24, -5.98, -5.975, -6.325, -6.35, -6.46, 
    -6.48, -6.93, -7.535, -7.795, -8.035, -8.045, -7.93, -8.735, -8.93, 
    -7.295, -6.155, -6.31, -5.095, -4.445, -5.165, -6.095, -5.32, -6.735, 
    -8.38, -9.31, -9.57, -9.25, -9.895, -9.365, -8.545, -8.21, -7.295, -6.67, 
    -7.195, -6.61, -6.67, -6.725, -6.145, -5.555, -5.355, -4.36, -3.695, 
    -4.14, -4.485, -4.5, -4.57, -4.555, -4.615, -4.52, -4.37, -4.4, -4.33, 
    -4.315, -4.195, -4.16, -4.23, -4.41, -4.47, -4.605, -4.95, -5.225, -4.84, 
    -4, -3.795, -2.98, -1.985, -2.375, -2.63, -2.42, -2.535, -4.08, -6.485, 
    -6.71, -5.935, -6.07, -6.475, -6.465, -6.67, -6.925, -7.095, -7.7, -7.6, 
    -7.435, -7.48, -7.89, -8.11, -8.09, -8, -7.58, -7.225, -6.825, -6.825, 
    -6.71, -6.68, -7.045, -8.085, -8.965, -9.575, -9.685, -9.85, -10.19, 
    -10.47, -11.075, -11.385, -11.22, -12.165, -12.885, -14.19, -14.465, 
    -13.165, -6.15, -5.99, -6.675, -5.78, -4.725, -6.39, -7.43, -8.135, 
    -8.98, -10.35, -10.75, -11.035, -12.695, -13.41, -13.825, -14.255, 
    -14.295, -14.6, -15.105, -13.685, -12.32, -11.06, -11.32, -10.655, -9.62, 
    -9.305, -8.37, -8.195, -6.635, -8.045, -7.84, -7.43, -8.675, -11.25, 
    -13.195, -11.835, -12.225, -12.505, -11.32, -11.215, -10.7, -10.465, 
    -10.26, -9.855, -9.795, -9.725, -9.865, -9.715, -8.72, -8.1, -7.4, -6.72, 
    -6.94, -8.03, -7.95, -7.94, -8.505, -8.735, -8.84, -8.865, -9.165, -9.31, 
    -9.26, -9.06, -9.1, -9.045, -8.615, -8.56, -8.64, -8.805, -8.88, -8.76, 
    -8.4, -7.845, -7.49, -7.125, -7.01, -6.955, -6.95, -6.745, -6.995, -7.18, 
    -7.28, -7.07, -7.095, -7.025, -6.625, -6.395, -6.305, -6.3, -6.215, 
    -6.22, -6.33, -6.355, -6.22, -5.985, -5.475, -5.3, -5.195, -4.985, -4.92, 
    -4.855, -5.115, -5.4, -5.455, -5.76, -5.695, -5.47, -5.305, -5.165, 
    -5.085, -5.23, -5.325, -5.285, -5.295, -5.315, -5.375, -5.275, -5.255, 
    -5.175, -4.885, -4.745, -4.825, -4.745, -4.745, -4.535, -5.295, -5.79, 
    -6.865, -8.16, -8.745, -9.715, -10.79, -9.655, -10.88,
  -7.355, -7.545, -6.75, -6.6, -6.515, -6.545, -7.34, -7.17, -5.715, -3.385, 
    -2.5, -2.31, -2.12, -1.97, -1.89, -2.04, -2.135, -3.33, -4.08, -4.8, 
    -5.035, -5.04, -4.9, -5.815, -5.1, -5.15, -5.315, -5.8, -6.785, -6.35, 
    -5.995, -4.845, -0.33, 1.05, 2.065, 2.82, 3.24, 4.18, 5.065, 4.925, 
    3.445, 2.475, 0.415, -2.325, -2.92, -3.28, -3.53, -2.68, -1.465, -2.74, 
    -1.81, -1.145, -0.18, -0.495, -0.52, 0.235, 1.205, 2.535, 2.73, 3.665, 
    4.295, 4.175, 4.94, 4.9, 4.45, 4.64, 2.975, 2.725, 2.615, 2.685, 2.435, 
    1.81, 0.91, 0.205, -0.235, -0.47, -0.515, -0.64, -0.845, -1.78, -2.05, 
    -1.92, -2.125, -1.23, -1.25, -1.145, -1.6, -1.23, -1.585, -1.585, -2.3, 
    -3.15, -3.33, -3.36, -3.455, -3.855, -4.075, -4.75, -4.96, -5.165, 
    -5.515, -5.835, -6.545, -6.57, -5.72, -5.005, -4.595, -4.815, -3.385, 
    -3.49, -4.83, -4.685, -4.665, -4.815, -4.99, -5.62, -5.855, -6.195, 
    -6.57, -7.72, -6.98, -8.075, -8.33, -7.45, -7.99, -9.205, -9.06, -7.505, 
    -3.675, -0.52, -1.075, 0.005, 0.47, 0.59, 1.325, 1.63, 1.59, -0.02, 
    -1.915, -3.25, -3.25, -2.425, -4.04, -5.65, -5.835, -5.745, -5.095, 
    -5.94, -6.22, -4.83, -5.01, -4.02, 1.03, 3.93, 4.6, 4.285, 5.385, 5.39, 
    5.855, 5.045, 3.88, 2.25, -0.07, -1.25, -1.275, -1.83, -2.23, -2.965, 
    -3.6, -4.115, -3.435, -3.18, -3.76, -4.225, -3.655, -3.03, -2.51, -2.165, 
    0.25, 0.005, 0.1, -0.37, -0.09, 0.575, -0.515, -1.49, -1.795, -1.965, 
    -2.835, -2.945, -2.88, -3.1, -3.305, -3.18, -3.02, -3.015, -2.87, -2.635, 
    -2.615, -2.5, -2.25, -1.475, -1.045, -0.975, -0.885, -0.44, 0.04, 0.575, 
    0.585, 0.22, -0.6, -1.41, -1.905, -2.355, -2.885, -3.295, -3.56, -3.7, 
    -3.8, -4.255, -4.765, -5.17, -5.03, -5.185, -4.64, -3.875, -3.515, 
    -1.445, -0.825, -1.09, -1.695, -2.995, -3.1, -3.2, -3.325, -3.35, -3.39, 
    -3.75, -3.445, -3.285, -3.715, -4.055, -3.645, -3.545, -3.24, -2.81, 
    -2.575, -2.42, -2.11, -1.765, -1.535, -1.51, -1.54, -1.775, -1.7, -0.625, 
    -0.39, -0.87, -1.65, -2.055, -2.42, -2.41, -2.55, -2.84, -2.545, -2.04, 
    -2.205, -2.17, -2.405, -3.215, -3.525, -3.61, 0.655, 3.6, 5.785, 6.57, 
    6.995, 7.15, 7.53, 7.385, 5.8, 4.335, 4.11, 4.4, 4.24, 4.335, 4.73, 
    4.535, 2.89, 1.555, 0.325, 0.35, 0.845, 0.995, 0.935, 1.355, 1.905, 
    4.155, 4.245, 4.125, 6.345, 5.6, 5.915, 5.98, 5.43, 4.75, 4.135, 3.435, 
    1.83, 1.76, 2.32, 1.64, 0.425, 0.01, -0.145, -0.32, -0.23, -0.18, -0.03, 
    0.285, 0.6, 1.02, 1.555, 2.43, 3, 4.035, 3.705, 3.68, 3.845, 3.64, 2.905, 
    3.01, 3.07, 3.265, 3.21, 2.86, 2.855, 2.865, 2.67, 2.83, 2.345, 1.865, 
    1.64, 1.73, 3.605, 3.61, 3.465, 3.61, 4.065, 4.53, 5.265, 5.195, 5.21, 
    4.105, 3.33, 3.12, 2.525, 1.895, 0.15, 1.09, 0, -0.015, -0.63, 0.365, 
    0.835, -0.315, -0.39, -0.23, 4.315, 6.37, 6.895, 7.54, 8.86, 9.645, 
    9.965, 10.18, 9.68, 7.155, 4.065, 3.22, 3.015, 2.745, 2.37, 2.38, 2.035, 
    2.295, 1.67, 3.37, 4.295, 3.935, 3.145, 3.32, 8.21, 11.115, 11.675, 
    12.655, 13.19, 13.435, 13.86, 13.49, 12.665, 10.17, 7.065, 5.96, 5.635, 
    5.365, 5.86, 5.51, 6.28, 7.3, 6.65, 6.65, 6.48, 6.695, 5.76, 5.82, 10.15, 
    11.875, 13.14, 14.395, 14.8, 14.755, 14.34, 14.805, 13.355, 10.935, 
    8.645, 7.925, 8.335, 8.8, 9.5, 9.395, 9.405, 9.295, 9.275, 8.95, 8.11, 
    6.99, 5.58, 2.68, 3.73, 6.09, 8.08, 7.55, 8.205, 8.445, 7.735, 7.105, 
    3.555, 1.365, 1.605, 0.555, -0.095, -0.245, -0.26, -0.435, -0.365, 
    -0.355, -0.08, -0.255, -0.205, -0.09, -0.065, -0.125, -0.135, 0.01, 
    1.385, 1.325, 2.04, 1.44, 0.56, 1.59, 2, 0.745, -0.065, -1.02, -1.85, 
    -2.13, -2.685, -2.695, -2.875, -2.955, -3.25, -3.665, -3.755, -3.6, 
    -3.76, -3.7, -0.905, -0.065, 1.235, 1.45, 1.37, 1.02, 2.045, 3.05, 2.44, 
    0.715, 0.185, -0.005, -0.605, -0.89, -0.365, -0.47, -0.855, -0.65, 
    -0.475, -0.29, -0.12, -0.145, -1.565, -1.24, -0.695, 0.885, 3.405, 3.905, 
    4.145, 5.08, 5.135, 4.29, 3.015, 1.875, 1.085, 0.55, 0.14, -0.35, -0.775, 
    -1.04, -1.3, -1.82, -2.17, -1.585, -2.265, -1.475, -1.1, -0.55, -0.065, 
    0.42, 1.105, 1.775, 1.865, 1.84, 1.32, 1.39, 1.325, 1.255, 0.875, 1.505, 
    1.655, 0.38, -0.1, -0.275, -0.385, -0.22, 0.45, 0.43, 0.49, 0.57, 0.58, 
    0.53, 0.44, 0.31, 0.385, 0.665, 1.135, 0.99, 1.275, 0.67, 0.04, -1.21, 
    -2.36, -3.435, -3.77, -4.13, -4.62, -4.36, -5.16, -5.175, -5.795, -6.895, 
    -7.15, -7.68, -8.83, -8.525, -5.37, -3.675, -2.575, -2.4, -1.495, -1.24, 
    -1.025, -0.9, -1.645, -3.29, -4.665, -5.31, -6.23, -6.83, -6.85, -6.555, 
    -6.935, -6.27, -5.78, -4.76, -4.385, -5.055, -4.825, -4.195, -2.995, 
    -0.53, 0.425, 0.46, 1.77, 2.12, 1.37, 1.625, 0.675, -0.295, -0.265, 0.47, 
    0.575, 0.845, 1.185, 2.2, 1.26, -1.705, -3.45, -4.61, -5.7, -7.2, -7.61, 
    -7.88, -8.115, -8.325, -8.22, -6.61, -5.275, -5.45, -5.67, -7.43, -8.115, 
    -9.05, -9.905, -9.425, -9.425, -9.975, -10.41, -10.37, -10.525, -10.585, 
    -10.59, -10.185, -10.37, -10.9, -10.375, -10.3, -9.47, -7.345, -4.955, 
    -4.905, -4.81, -3.835, -3.385, -4.11, -4.87, -6.115, -6.84, -7.425, 
    -7.925, -8.435, -8.58, -8.355, -8.895, -9.32, -10.21, -11.555, -10.74, 
    -9.74, -11.12, -11.795, -8.96, -8.105, -6.325, -5.97, -5.05, -4.475, 
    -5.55, -6.345, -7.165, -8.095, -8.82, -9.12, -9.48, -9.46, -9.425, 
    -9.385, -9.26, -8.82, -8.485, -8.135, -7.27, -6.12, -5.78, -4.615, 
    -3.995, -4.02, -4.47, -3.84, -3.655, -3.445, -2.9, -2.355, -2.185, 
    -2.095, -1.985, -1.8, -1.595, -1.53, -1.515, -1.49, -1.565, -1.435, 
    -1.435, -1.68, -1.955, -2.365, -2.435, -2.37, -1.365, -0.055, 0.575, 1.5, 
    3.035, 3.68, 4.335, 4.95, 3.63, 1.775, 0.865, 0.36, 0.275, 0.995, 1.82, 
    1.785, 1.4, 1.36, 1.285, 1.6, 1.835, 1.875, 1.515, 1.73, 3.245, 4.875, 
    5.565, 6.04, 5.82, 5.32, 5.02, 4.055, 4.01, 3.235, 2.145, 1.935, 1.62, 
    1.66, 1.345, 1.35, 0.745, 0.8, 0.725, 0.695, 0.09, 0.1, -0.44, -0.665, 
    1.735, 4.885, 5.61, 6.485, 6.69, 6.055, 6.27, 5.845, 5.125, 3.245, 1.01, 
    0.41, 1.095, 0.325, 0.5, 0.305, 0.655, 1.325, 1.02, 1.255, 0.355, 0.56, 
    0.72, 0.96, 3.15, 5.19, 5.59, 7.01, 7.335, 7.925, 7.875, 7.895, 6.835, 
    4.98, 2.54, 0.655, 0.6, 0.4, 0.27, 0.49, 0.76, 0.82, 1.415, 3.575, 4.175, 
    1.61, 1.81, 1.805, 5.895, 10.93, 11.875, 12.64, 13.65, 14.125, 14.33, 
    13.455, 11.69, 8.375, 6.52, 6.475, 8.25, 8.96, 7.66, 7.7, 7.52, 7.625, 
    7.815, 6.98, 4.965, 3.055, 2.155, 4.905, 7.49, 9.84, 11.135, 12.03, 
    12.36, 11.785, 12.515, 10.92, 10.01, 8.255, 7.295, 6.835, 7.165, 7.89, 
    8.21, 7.47, 6.67, 6.075, 6.055, 5.65, 5.05, 4.79, 4.53, 4.405, 4.635, 
    6.24, 6.61, 6.805, 7.015, 6.83, 6.02, 4.875, 4.105, 3.2, 2.305, 2.36, 
    2.155, 1.6, 1.145, 0.875, 0.415, -0.01, -0.35, -0.21, -0.37, -0.445, 
    -0.4, -0.04, 0.475, 2.315, 3.425, 4.885, 5.01, 3.305, 2.65, 1.91, 2.11, 
    1.01, -0.785, -2.23, -2.46, -2.97, -3.2, -2.71, -2.51, -2.93, -3.775, 
    -4.095, -4.535, -4.84, -6.07, -6.715, -3.515, -0.39, -0.05, -0.225, 0.32, 
    0.97, 1.155, 0.89, 0.04, -2.045, -3.91, -4.535, -4.6, -5.05, -5.16, 
    -4.72, -4.505, -5.255, -6.435, -6.42, -5.605, -5.01, -5.03, -4.77, 
    -2.195, 2.48, 4.08, 5.16, 5.565, 5.865, 6.11, 5.7, 4.06, 1.125, 0.435, 
    1.28, 0.965, 0.3, 1.215, 0.53, 0.51, 1.36, 0.055, -0.23, -0.62, 0, 0.895, 
    0.905, 1.045, 2.225, 3.185, 4.6, 4.88, 5.415, 4.655, 4.425, 3.8, 1.905, 
    -0.445, -1.38, -1.93, -1.92, 0.985, 2.22, 2.435, 1.735, 1.81, 2.32, 
    2.415, 1.915, 0.91, 2.285, 2.85, 5.575, 7.23, 8.69, 8.46, 7.6, 6.61, 6.31, 
    6.02, 5.235, 4.925, 4.94, 4.37, 3.765, 5.105, 5.15, 4.895, 4.455, 3.955, 
    3.905, 3.905, 3.665, 3.23, 2.34, 2.375, 2.05, 0.97, 0.635, -1.855, -2.95, 
    -3.085, -3.63, -4.23, -5.015, -5.825, -6.425, -7.33, -8.405, -8.91, 
    -8.615, -9.645, -10.04, -10.88, -11.45, -11.965, -12.235, -12.515, 
    -12.415, -10.93, -8.25, -6.695, -6.955, -5.96, -7.365, -6.795, -7.075, 
    -7.945, -9.305, -11.035, -11.44, -11.825, -11.58, -12.035, -12.755, 
    -12.61, -11.075, -10.5, -10.245, -9.655, -9.535, -9.825, -9.65, -9.095, 
    -8.31, -7.095, -7.035, -6.855, -7.495, -8.515, -9.36, -9.965, -10.825, 
    -11.33, -11.56, -11.925, -12.32, -12.825, -12.88, -13.815, -14.32, 
    -14.955, -14.53, -14.415, -14.87, -14.375, -14.77, -14.145, -10.085, 
    -9.09, -8.33, -6.735, -7.955, -7.56, -8.015, -9.275, -10.56, -12.09, 
    -12.675, -13.005, -12.425, -11.535, -10.825, -10.895, -10.755, -10.785, 
    -10.695, -10.23, -10.43, -10.04, -9.725, -7.485, -1.285, -0.29, -0.16, 
    -0.38, -0.045, -0.255, 0.37, -1.49, -2.965, -3.435, -3.87, -3.155, 
    -2.305, -2.33, -2.59, -2.8, -1.925, -1.735, -1.4, -2.195, -2.29, -0.96, 
    -2.005, 0.03, 5.11, 6.15, 6.175, 7.57, 7.14, 7.885, 6.83, 4.14, 0.645, 
    -0.96, -0.375, -0.04, -0.23, -0.145, -0.28, -1.02, 0.615, 0.77, 0.62, 
    0.16, 0.315, -0.91, -2.27, -0.615, 4.14, 4.54, 3.83, 3.195, 3.43, 3.36, 
    2.745, 0.845, -0.315, -1.91, -2.33, -2.745, -3.535, -4.07, -5.01, -5.47, 
    -5.905, -7.04, -7.385, -7.685, -7.2, -6.375, -6.535, -5.69, -3.28, 
    -0.525, 0.79, 0.905, 1.02, 1.56, 1.49, -0.495, -2.175, -2.895, -3.095, 
    -3.4, -2.645, -1.965, -2.055, -2.165, -2.97, -4.335, -3.815, -2.18, 0.21, 
    0.665, 0.43, 0.655, 3.58, 3.495, 4.245, 4.465, 4.85, 4.59, 4.26, 3.67, 
    2.045, 1.785, 2.055, 2.625, 2.445, 2.395, 2.105, 1.475, 0.92, -0.795, 
    -2.14, -3.39, -5.35, -5.66, -5.84, -6.37, -6.355, -6.04, -6.16, -6.745, 
    -6.245, -6.955, -7.37, -8, -8.72, -9.125, -9.62, -10.505, -11.24, -11.81, 
    -12.43, -12.6, -13.06, -13.38, -11.865, -10.825, -10.53, -11.27, -10.905, 
    -9.55, -7.595, -4.085, -3.155, -4.43, -5.375, -6.38, -6.51, -6.2, -7.65, 
    -8.285, -8.77, -9.165, -9.735, -10.02, -10.195, -10.51, -10.71, -10.93, 
    -11.065, -11, -11.06, -11.17, -11.32, -11.375, -10.61, -9.92, -8.895, 
    -8.965, -8.75, -8.755, -9.17, -10.595, -10.675, -10.62, -11.175, -11.345, 
    -11.39, -11.695, -11.66, -11.335, -11.495, -12.24, -12.115, -12.18, 
    -12.14, -11.995, -11.935, -10.885, -7.475, -4.39, -2.31, -2.73, -2.565, 
    -1.045, -1.31, -3.53, -4.64, -4.62, -4.335, -5.515, -5.86, -5.425, 
    -5.865, -5.865, -5.38, -5.42, -5.465, -5.11, -4.655, -5, -5.305, -3.68, 
    0.3, 1.87, 2.7, 3.505, 3.69, 4.08, 3.49, 1.735, -0.97, -2.08, -2.675, 
    -3.06, -3.27, -3.89, -3.07, -1.875, -2.305, -2.15, -2.1, -2.715, -2.985, 
    -0.955, -0.215, 0.515, 5.195, 8.785, 9.225, 8.35, 8.725, 7.705, 6.05, 
    3.71, 0.975, -1.16, -2.095, -1.58, -1.835, -0.91, -0.03, -1.605, -1.17, 
    -1.895, -1.175, -1.545, -2.025, -3.73, -3.86, -3.345, 2.315, 3.785, 
    5.015, 4.19, 3.585, 3.145, 2.52, 1.955, -1.575, -3.39, -3.575, -3.205, 
    -2.665, -2.745, -2.525, -2.835, -2.58, -2.665, -2.57, -3.01, -3.335, 
    -3.565, -3.855, -3.535, -2.955, -1.765, 0.75, 1.5, 1.08, 0.455, 0.315, 
    -1.165, -2.665, -3.43, -4.005, -4.715, -5.455, -5.78, -6.79, -7.465, 
    -7.335, -7.735, -7.89, -6.925, -6.36, -5.835, -6.605, -6.105, -2.23, 
    -0.71, 0.665, 1.175, 1.4, 1.33, 0.61, -1.795, -3.185, -4.505, -5.175, 
    -5.71, -6.015, -5.5, -5.5, -5.585, -5.24, -4.56, -4.76, -4.69, -4.35, 
    -4.465, -4.26, -3.565, 1.83, 3.505, 2.76, 2.385, 2.26, 2.495, 1.51, 
    0.325, -1.195, -1.64, -2.145, -2.565, -3.025, -3.54, -3.24, -3.705, 
    -4.01, -4.6, -4.815, -4.81, -4.86, -5.15, -5.755, -5.32, -3.705, -2.425, 
    -1.77, -2.05, -3.41, -4.075, -4.72, -5.075, -5.605, -6.04, -6.7, -7.5, 
    -7.795, -8.12, -8.675, -10.235, -11.22, -11.485, -12.015, -12.63, -13.78, 
    -15.085, -15.58, -14.845, -11.125, -8.695, -6.685, -6.2, -6.495, -6.385, 
    -7.42, -9.66, -11.865, -13.28, -14.14, -14.65, -15.61, -16.54, -16.78, 
    -17.69, -17.96, -18.28, -18.675, -19.345, -19.56, -19.125, -19.805, 
    -19.305, -14.49, -11.81, -11.34, -11.38, -10.775, -10.575, -10.95, 
    -12.405, -14.26, -15.32, -16.83, -15.885, -16.525, -16.755, -16.51, 
    -15.7, -15.335, -15.35, -15.14, -14.785, -14.17, -13.585, -13.835, 
    -14.24, -12.725, -10.805, -9.535, -7.9, -7.18, -6.33, -7.795, -9.215, 
    -10.115, -9.975, -9.47, -9.36, -9.225, -8.995, -9.485, -9.485, -9.63, 
    -10.185, -11.245, -9.905, -9.77, -10.84, -12.165, -12.645, -12.71, 
    -12.485, -11.98, -10.905, -10.755, -11.565, -12.84, -14.165, -15.435, 
    -15.755, -15.655, -16.355, -17.17, -16.77, -16.02, -15.865, -16.38, 
    -17.825, -18.595, -19.02, -19.315, -19.555, -19.755, -19.985, -19.705, 
    -19.19, -18.81, -18.725, -18.26, -18.495, -18.97, -19.66, -20.705, 
    -21.335, -21.745, -22.295, -23.25, -24.245, -24.665, -24.505, -24.485, 
    -24.37, -24.205, -23.345, -22.25, -22.24, -22.17, -22.07, -21.72, 
    -18.895, -19.35, -17.555, -14.885, -12.675, -15.025, -18.625, -17.785, 
    -16.245, -17.095, -16.09, -16.875, -17.51, -18.045, -18.28, -18.3, 
    -18.415, -17.535, -16.975, -17.025, -17.1, -17.755, -18.285, -18.105, 
    -18.125, -17.525, -17.12, -17.48, -18.1, -18.54, -19.775, -20.585, 
    -21.17, -21.385, -21.095, -21.08, -21.235, -20.99, -20.805, -20.515, 
    -20.42, -20.185, -20.075, -20.405, -20.71, -21.015, -20.97, -20.575, 
    -20.225, -19.76, -19.475, -19.22, -19.465, -19.27, -19.115, -19.405, 
    -19.44, -19.37, -19.37, -19.395, -19.415, -19.415, -19.275, -19.17, 
    -19.21, -19.08, -18.99, -18.95, -18.815, -19.28, -18.905, -15.135, 
    -12.275, -11.595, -10.325, -10.455, -11.855, -12.435, -14.485, -15.87, 
    -17.055, -16.975, -16.375, -16.115, -16.07, -16, -15.48, -15.11, -14.535, 
    -14.875, -14.745, -14.215, -13.755, -13.425, -12.825, -10.51, -7.39, 
    -5.575, -4.445, -4.69, -4.975, -6.65, -7.895, -9.725, -11.065, -10.655, 
    -11.37, -10.1, -9.975, -9.885, -9.42, -9.41, -8.945, -8.61, -8.47, 
    -8.175, -7.835, -7.43, -7.385, -7.315, -6.92, -6.52, -6.23, -5.77, -5.79, 
    -6.225, -6.285, -6.125, -5.98, -5.755, -5.645, -5.51, -5.42, -5.425, 
    -5.535, -5.615, -5.5, -5.315, -5.195, -5.08, -5.12, -5.225, -5.365, 
    -5.59, -5.365, -5.44, -5.41, -5.505, -5.91, -6.135, -6.27, -6.38, -6.515, 
    -6.58, -6.55, -6.56, -6.645, -6.965, -7.265, -7.38, -7.825, -7.89, -7.78, 
    -7.7, -7.755, -7.95, -8.075, -8.12, -8.325, -8.255, -7.81, -8.43, -8.73, 
    -8.65, -9.255, -9.505, -9.465, -9.515, -9.92, -10.06, -10.07, -10.025, 
    -9.935, -9.81, -9.62, -8.785, -8.325, -8.485, -8.735, -8.785, -8.92, 
    -5.815, -4.445, -2.155, -2.13, -4.205, -4.08, -5.545, -6.225, -6.72, 
    -6.51, -6.09, -5.84, -5.775, -5.79, -5.185, -5.145, -4.935, -4.48, -4.06, 
    -3.765, -3.84, -4.545, -4.635, -3.765, -2.795, -2.095, -2.21, -2.855, 
    -3.545, -3.3, -3.06, -2.925, -3.525, -3.695, -3.95, -3.685, -3.495, 
    -3.18, -2.925, -3.41, -3.555, -3.325, -3.215, -3.42, -3.67, -3.945, 
    -4.09, -4.305, -4.125, -3.16, -3.65, -3.36, -2.73, -2.61, -3.21, -4.645, 
    -5.35, -5.675, -5.55, -5.51, -5.575, -5.635, -6.055, -6.94, -7.69, 
    -8.405, -9.185, -8.205, -7.705, -7.895, -7.725, -7.58, -6.49, -3.005, 
    -4.335, -3.93, -4.2, -3.965, -5.115, -6.095, -7.21, -7.88, -8.145, 
    -8.285, -8.885, -8.875, -8.96, -9.115, -8.93, -9.305, -9.47, -9.33, 
    -7.835, -7.315, -7.565, -7.18, -6.55, -5.3, -4.76, -4.48, -4.66, -4.61, 
    -4.58, -4.835, -5.255, -5.445, -5.325, -5.35, -5.245, -5.005, -4.79, 
    -4.74, -4.655, -4.06, -3.845, -3.125, -3.29, -2.995, -3.185, -3.31, 
    -2.025, 1.175, 2.505, 3.175, 3.145, 2.57, 1.095, -1.35, -2.875, -3.63, 
    -4.415, -5.305, -5.74, -4.94, -4.63, -4.425, -4.875, -5.035, -4.79, 
    -5.865, -5.805, -5.955, -5.34, -5.38, -2.91, -0.385, -0.27, 0.215, -0.42, 
    -0.215, -1.255, -2.87, -4.465, -5.465, -7.125, -7.495, -6.945, -5.57, 
    -5.24, -4.35, -4.25, -4.575, -4.62, -4.525, -4.58, -5.09, -5.075, -5.31, 
    -5.065, -4.22, -4.815, -5.265, -5.525, -6.25, -6.02, -6.115, -6.55, 
    -6.92, -6.215, -5.89, -5.82, -5.755, -5.795, -6.735, -8.43, -9.43, -8.76, 
    -8.13, -7.59, -7.745, -8.195, -8.035, -7.89, -7.93, -8.515, -8.45, -8.89, 
    -9.35, -10.29, -11.62, -12.92, -13.94, -14.675, -15.21, -16, -16.61, 
    -16.38, -17.19, -17.32, -17.855, -17.57, -18.915, -18.505, -17.815, 
    -18.93, -19.07, -15.53, -13.015, -12.67, -12.56, -12.655, -11.455, 
    -12.965, -14.29, -15.45, -15.815, -15.785, -15.355, -14.63, -14.145, 
    -14.09, -14.285, -14.1, -13.745, -13.875, -14.36, -14.435, -13.25, -12.4, 
    -12.58, -11.29, -8.965, -8.625, -8.975, -9.55, -10.125, -11.08, -11.315, 
    -12.695, -13.315, -13.875, -13.795, -14.37, -14.84, -13.87, -13.465, 
    -13.915, -14.755, -15.205, -15.305, -15.57, -15.355, -15.43, -14.65, 
    -9.12, -4.545, -3, -5.655, -6.365, -6.82, -6.97, -8.125, -10.44, -12.505, 
    -12.785, -12.57, -11.98, -11.945, -12.24, -11.8, -11.285, -10.035, 
    -10.09, -9.615, -10.11, -10.335, -9.92, -10.165, -7.91, -5.725, -5.41, 
    -5.31, -5.18, -5.97, -6.53, -7.595, -8.935, -9.815, -10.375, -10.545, 
    -11.495, -11.895, -12.705, -12.995, -12.85, -13.365, -12.865, -13.145, 
    -13.335, -13.625, -11.99, -12.155, -7.805, -2.85, -2.62, -2.51, -2.495, 
    -2.89, -3.86, -5.75, -8.58, -10.49, -9.89, -9.2, -9.57, -9.025, -9.41, 
    -9.21, -10.37, -10.85, -10.56, -9.405, -9.39, -10.125, -10.545, -9.535, 
    -8.555, -7.765, -8.935, -8.975, -8.225, -8.225, -8.305, -9.36, -10.3, 
    -10.46, -10.32, -10.325, -10.44, -10.57, -10.73, -10.81, -10.83, -10.85, 
    -10.68, -10.515, -10.485, -10.46, -10.375, -10.2, -9.87, -9.71, -9.97, 
    -10.115, -10.29, -10.265, -10.525, -10.655, -10.83, -11.13, -11.32, 
    -11.45, -11.365, -11.41, -11.175, -11, -11.05, -11.16, -11.21, -11.25, 
    -11.325, -11.46, -11.74, -11.78, -11.23, -10.245, -9.775, -9.115, -8.925, 
    -10.265, -10.64, -11.025, -11.22, -11.205, -11.165, -11, -10.64, -10.21, 
    -9.67, -8.725, -7.44, -7.26, -7.165, -6.45, -6.07, -5.98, -5.965, -5.635, 
    -4.63, -3.835, -3.85, -3.82, -4.06, -3.585, -4.02, -4.765, -5.095, -5.26, 
    -5.36, -5, -4.545, -4.355, -4.075, -4.35, -4.48, -4.435, -4.39, -4.57, 
    -4.73, -5.175, -5.51, -6.235, -6.595, -6.35, -6.12, -6.375, -5.735, 
    -6.26, -6.19, -6.82, -7.175, -7.385, -7.775, -8.295, -8.16, -8.425, 
    -8.16, -7.82, -7.76, -7.835, -7.975, -8.065, -8.135, -8.09, -7.875, 
    -7.91, -7.56, -6.925, -5.675, -5.265, -4.71, -4.275, -5.165, -7.075, 
    -7.53, -8.385, -10.07, -11.04, -9.97, -9.465, -9.525, -9.72, -9.175, 
    -8.805, -9.18, -8.68, -9.065, -9.46, -9.745, -8.465, -6.73, -3.945, 
    -0.485, -0.495, -0.645, -2.17, -4.61, -5.76, -6.04, -6.25, -6.28, -5.96, 
    -6.185, -5.615, -5.485, -5.62, -5.33, -5.25, -5.07, -4.695, -4.665, 
    -4.62, -4.345, -4.385, -4.2, -4.09, -4.535, -3.27, -3.08, -3.26, -3.99, 
    -4.615, -5.075, -5.045, -4.375, -4.35, -4.355, -4.49, -4.785, -4.645, 
    -4.725, -4.53, -4.265, -4.075, -3.99, -3.95, -3.695, -3.64, -3.775, 
    -3.84, -3.81, -3.76, -3.865, -4.39, -4.74, -5.52, -6.44, -7.42, -7.99, 
    -8.725, -10.68, -12.035, -12.77, -12.49, -13.635, -15.155, -15.77, 
    -16.06, -16.15, -15.66, -15.92, -15.74, -12.88, -9.905, -6.055, -4.78, 
    -5.285, -5.765, -7.07, -8.32, -10.375, -12.445, -12.86, -12.95, -13.015, 
    -12.6, -12.31, -11.595, -11.38, -11.495, -11.11, -11.01, -10.505, -10.46, 
    -10.64, -10.375, -7.355, -3.06, -0.025, 0.585, -1.085, -1.615, -2.14, 
    -2.935, -4.09, -4.345, -5.01, -4.615, -4.715, -4.73, -4.525, -4.585, 
    -4.71, -5.085, -4.83, -4.06, -4.135, -4.375, -4.645, -5.415, -4.645, 
    -2.545, -1.125, -0.895, -0.94, -1.635, -2.395, -2.705, -3.54, -4.98, 
    -4.475, -4.38, -4.09, -5.535, -5.845, -5.85, -4.81, -4.02, -4.13, -4.63, 
    -5.645, -5.195, -5.64, -5.865, -2.765, 0.66, 1.53, 1.22, 1.9, 1.68, 1.07, 
    -0.37, -1.655, -3.4, -4.36, -4.665, -4.765, -4.8, -4.94, -5.55, -5.315, 
    -5.13, -4.915, -5.165, -5.695, -5.65, -5.645, -5.63, -1.34, 2.43, 3.78, 
    4.19, 3.38, 3.8, 3.395, 1.47, 0.345, -0.085, -0.675, -0.12, -2.305, 
    -4.25, -4.78, -4.225, -4.34, -5.215, -5.575, -2.12, -3.445, -1.35, 
    -0.435, -0.095, 1.43, 1.76, 2.09, 2.54, 2.19, 1.905, 1.185, 1.175, 
    -0.655, -1.435, -2.045, -1.88, -3.135, -3.9, -3.785, -2.76, -2.755, 
    -2.575, -3.11, -4.3, -5.945, -6.455, -6.14, -5.77, -3.155, 0.405, 2.715, 
    2.23, 2.61, 0.42, 1.26, -0.115, -1.685, -2.155, -2.805, -3.24, -3.125, 
    -3.45, -4.3, -4.965, -5.03, -5.665, -5.7, -5.585, -5.795, -5.925, -6.055, 
    -6.155, -5.78, -5.09, -5.12, -4.5, -4.32, -4.195, -4.57, -5.32, -6.03, 
    -6.63, -7.41, -8.055, -8.335, -8.65, -8.58, -8.6, -9.29, -10.37, -10.12, 
    -9.49, -8.435, -8.325, -9.545, -7.535, -6.17, -4.84, -3.28, -2.545, 
    -2.07, -1.18, -1.835, -2.55, -2.56, -2.47, -2.72, -2.68, -3.175, -3.03, 
    -2.35, -2.535, -3.365, -3.07, -3.2, -3.105, -4.345, -3.715, -3.79, 
    -3.585, -1.015, 0.52, 2.87, 3.41, 2.845, 1.565, 1.67, 0.03, -2.025, 
    -2.87, -3.785, -3.61, -3.735, -3.275, -2.905, -3.425, -2.73, -3.705, 
    -3.81, -4.375, -5.085, -6.665, -5.465, -4.25, -1.75, 1.065, 0.805, 1.4, 
    2.235, 2.115, 1.685, -0.19, -2.595, -4.095, -4.015, -3.665, -3.205, 
    -3.03, -2.985, -3.485, -4.155, -4.565, -5.53, -5.695, -4.95, -5.59, 
    -5.92, -5.84, -5.445, -4.705, -4.615, -3.24, -3.86, -3.725, -4.13, -4.04, 
    -4.295, -4.435, -4.19, -4.33, -4.815, -5.005, -5.065, -4.825, -4.8, 
    -4.64, -4.24, -4.485, -4.825, -4.995, -5.245, -5.265, -5.22, -5.775, 
    -5.79, -5.325, -4.55, -5.65, -5.77, -5.91, -7.145, -7.855, -9.365, -8.31, 
    -7.795, -7.275, -7.145, -7.52, -7.775, -7.36, -7.85, -8.25, -8.15, -8.14, 
    -8.6, -8.595, -7.36, -5.85, -4.705, -5.065, -5.045, -5.975, -5.795, 
    -5.55, -6.68, -7.605, -8.11, -7.86, -7.685, -7.485, -7.135, -7.315, 
    -7.36, -7.205, -6.965, -6.82, -6.835, -6.99, -6.895, -6.84, -6.525, 
    -6.02, -5.675, -4.24, -4.675, -4.665, -4.695, -5.27, -6.405, -7.235, 
    -7.1, -7.345, -7.725, -7.48, -7.275, -7.79, -7.68, -7.6, -7.385, -6.56, 
    -5.955, -6.11, -6.545, -6.635, -6.515, -6.17, -5.305, -5.655, -6.005, 
    -6.695, -7.035, -7.16, -7.205, -7.37, -7.59, -7.7, -7.82, -8.26, -8.495, 
    -8.565, -8.605, -8.81, -9.19, -9.41, -9.475, -9.51, -9.555, -9.64, -9.5, 
    -9.35, -9.2, -9.22, -9.44, -9.615, -9.78, -9.78, -9.685, -9.65, -9.625, 
    -9.6, -9.625, -9.74, -9.875, -9.965, -10.075, -10.175, -10.23, -10.215, 
    -10.255, -10.31, -10.31, -10.375, -10.22, -9.755, -8.63, -7.215, -8.505, 
    -9.28, -9.46, -10.105, -10.5, -10.91, -11.29, -11.585, -11.655, -11.925, 
    -12.14, -12.165, -11.54, -11.055, -11.17, -11.26, -10.815, -10.49, 
    -10.505, -10.025, -9.39, -9.115, -8.83, -8.345, -6.725, -6.045, -5.165, 
    -5.88, -7.2, -7.63, -7.795, -8.485, -10.6, -11.19, -9.17, -8.75, -9.605, 
    -10.255, -10.735, -10.06, -8.325, -6.455, -6.355, -6.43, -5.34, -3.955, 
    -2.875, -3.755, -3.085, -2.67, -2.3, -3.165, -4.445, -5.105, -5.345, 
    -5.525, -6.06, -6.5, -7.16, -7.35, -7.11, -8.16, -8.68, -8.495, -8.6, 
    -8.165, -7.945, -8.435, -6.715, -4.175, -2.98, -2.245, -2.635, -2.99, 
    -3.59, -4.015, -5.26, -6.64, -6.955, -6.945, -6.925, -6.8, -7.245, -7.65, 
    -8, -8.105, -8.07, -7.99, -8.055, -8.935, -9.44, -9.425, -6.345, -4.485, 
    -3.795, -3.12, -2.88, -2.25, -2.125, -3.3, -5.79, -7.66, -8.255, -8.985, 
    -9.48, -9.625, -10.43, -10.325, -9.5, -10.63, -10.7, -10.325, -10.52, 
    -10.815, -10.675, -10.165, -6.18, -3.14, -1.37, -1.145, -0.9, -0.62, 
    -0.66, -3.105, -4.88, -6.73, -6.945, -7.765, -8.805, -8.975, -8.825, 
    -8.2, -7.88, -9.39, -8.385, -8.9, -7.305, -7.37, -9.75, -9.985, -6.56, 
    -1.025, 1.22, 1.44, 0.785, 0.615, 0.5, -1.65, -3.605, -4.805, -5.71, 
    -5.435, -5.24, -5.53, -5.61, -5.725, -6.06, -6.46, -6.985, -7.275, 
    -7.265, -7.285, -7.25, -7.255, -7.085, -6.685, -6.695, -6.635, -6.77, 
    -6.92, -6.815, -7.225, -7.32, -7.365, -7.32, -7.345, -7.475, -7.72, 
    -7.725, -7.9, -8.01, -8.005, -8.005, -8.155, -8.295, -8.405, -8.615, 
    -8.675, -8.375, -7.33, -6.57, -6.145, -7.515, -6.66, -5.42, -6.335, 
    -7.645, -8.825, -9.915, -11.955, -11.91, -11.31, -10.255, -10.925, 
    -10.965, -10.295, -9.375, -9.245, -9.375, -9.755, -10.95, -10.68, -6.425, 
    -0.755, -0.125, -1.15, -2.785, -3.34, -3.385, -3.89, -4.725, -6.705, 
    -7.995, -7.465, -7.3, -7.64, -9.24, -9.84, -10.31, -9.99, -9.83, -9.6, 
    -9.3, -8.495, -7.625, -6.185, -4.885, -5.4, -4.21, -1.24, -1.065, -1.255, 
    -1.425, -2.215, -3.815, -5.24, -5.98, -5.975, -6.325, -6.35, -6.46, 
    -6.48, -6.93, -7.535, -7.795, -8.035, -8.045, -7.93, -8.735, -8.93, 
    -7.295, -6.155, -6.31, -5.095, -4.445, -5.165, -6.095, -5.32, -6.735, 
    -8.38, -9.31, -9.57, -9.25, -9.895, -9.365, -8.545, -8.21, -7.295, -6.67, 
    -7.195, -6.61, -6.67, -6.725, -6.145, -5.555, -5.355, -4.36, -3.695, 
    -4.14, -4.485, -4.5, -4.57, -4.555, -4.615, -4.52, -4.37, -4.4, -4.33, 
    -4.315, -4.195, -4.16, -4.23, -4.41, -4.47, -4.605, -4.95, -5.225, -4.84, 
    -4, -3.795, -2.98, -1.985, -2.375, -2.63, -2.42, -2.535, -4.08, -6.485, 
    -6.71, -5.935, -6.07, -6.475, -6.465, -6.67, -6.925, -7.095, -7.7, -7.6, 
    -7.435, -7.48, -7.89, -8.11, -8.09, -8, -7.58, -7.225, -6.825, -6.825, 
    -6.71, -6.68, -7.045, -8.085, -8.965, -9.575, -9.685, -9.85, -10.19, 
    -10.47, -11.075, -11.385, -11.22, -12.165, -12.885, -14.19, -14.465, 
    -13.165, -6.15, -5.99, -6.675, -5.78, -4.725, -6.39, -7.43, -8.135, 
    -8.98, -10.35, -10.75, -11.035, -12.695, -13.41, -13.825, -14.255, 
    -14.295, -14.6, -15.105, -13.685, -12.32, -11.06, -11.32, -10.655, -9.62, 
    -9.305, -8.37, -8.195, -6.635, -8.045, -7.84, -7.43, -8.675, -11.25, 
    -13.195, -11.835, -12.225, -12.505, -11.32, -11.215, -10.7, -10.465, 
    -10.26, -9.855, -9.795, -9.725, -9.865, -9.715, -8.72, -8.1, -7.4, -6.72, 
    -6.94, -8.03, -7.95, -7.94, -8.505, -8.735, -8.84, -8.865, -9.165, -9.31, 
    -9.26, -9.06, -9.1, -9.045, -8.615, -8.56, -8.64, -8.805, -8.88, -8.76, 
    -8.4, -7.845, -7.49, -7.125, -7.01, -6.955, -6.95, -6.745, -6.995, -7.18, 
    -7.28, -7.07, -7.095, -7.025, -6.625, -6.395, -6.305, -6.3, -6.215, 
    -6.22, -6.33, -6.355, -6.22, -5.985, -5.475, -5.3, -5.195, -4.985, -4.92, 
    -4.855, -5.115, -5.4, -5.455, -5.76, -5.695, -5.47, -5.305, -5.165, 
    -5.085, -5.23, -5.325, -5.285, -5.295, -5.315, -5.375, -5.275, -5.255, 
    -5.175, -4.885, -4.745, -4.825, -4.745, -4.745, -4.535, -5.295, -5.79, 
    -6.865, -8.16, -8.745, -9.715, -10.79, -9.655, -10.88,
  -7.355, -7.545, -6.75, -6.6, -6.515, -6.545, -7.34, -7.17, -5.715, -3.385, 
    -2.5, -2.31, -2.12, -1.97, -1.89, -2.04, -2.135, -3.33, -4.08, -4.8, 
    -5.035, -5.04, -4.9, -5.815, -5.1, -5.15, -5.315, -5.8, -6.785, -6.35, 
    -5.995, -4.845, -0.33, 1.05, 2.065, 2.82, 3.24, 4.18, 5.065, 4.925, 
    3.445, 2.475, 0.415, -2.325, -2.92, -3.28, -3.53, -2.68, -1.465, -2.74, 
    -1.81, -1.145, -0.18, -0.495, -0.52, 0.235, 1.205, 2.535, 2.73, 3.665, 
    4.295, 4.175, 4.94, 4.9, 4.45, 4.64, 2.975, 2.725, 2.615, 2.685, 2.435, 
    1.81, 0.91, 0.205, -0.235, -0.47, -0.515, -0.64, -0.845, -1.78, -2.05, 
    -1.92, -2.125, -1.23, -1.25, -1.145, -1.6, -1.23, -1.585, -1.585, -2.3, 
    -3.15, -3.33, -3.36, -3.455, -3.855, -4.075, -4.75, -4.96, -5.165, 
    -5.515, -5.835, -6.545, -6.57, -5.72, -5.005, -4.595, -4.815, -3.385, 
    -3.49, -4.83, -4.685, -4.665, -4.815, -4.99, -5.62, -5.855, -6.195, 
    -6.57, -7.72, -6.98, -8.075, -8.33, -7.45, -7.99, -9.205, -9.06, -7.505, 
    -3.675, -0.52, -1.075, 0.005, 0.47, 0.59, 1.325, 1.63, 1.59, -0.02, 
    -1.915, -3.25, -3.25, -2.425, -4.04, -5.65, -5.835, -5.745, -5.095, 
    -5.94, -6.22, -4.83, -5.01, -4.02, 1.03, 3.93, 4.6, 4.285, 5.385, 5.39, 
    5.855, 5.045, 3.88, 2.25, -0.07, -1.25, -1.275, -1.83, -2.23, -2.965, 
    -3.6, -4.115, -3.435, -3.18, -3.76, -4.225, -3.655, -3.03, -2.51, -2.165, 
    0.25, 0.005, 0.1, -0.37, -0.09, 0.575, -0.515, -1.49, -1.795, -1.965, 
    -2.835, -2.945, -2.88, -3.1, -3.305, -3.18, -3.02, -3.015, -2.87, -2.635, 
    -2.615, -2.5, -2.25, -1.475, -1.045, -0.975, -0.885, -0.44, 0.04, 0.575, 
    0.585, 0.22, -0.6, -1.41, -1.905, -2.355, -2.885, -3.295, -3.56, -3.7, 
    -3.8, -4.255, -4.765, -5.17, -5.03, -5.185, -4.64, -3.875, -3.515, 
    -1.445, -0.825, -1.09, -1.695, -2.995, -3.1, -3.2, -3.325, -3.35, -3.39, 
    -3.75, -3.445, -3.285, -3.715, -4.055, -3.645, -3.545, -3.24, -2.81, 
    -2.575, -2.42, -2.11, -1.765, -1.535, -1.51, -1.54, -1.775, -1.7, -0.625, 
    -0.39, -0.87, -1.65, -2.055, -2.42, -2.41, -2.55, -2.84, -2.545, -2.04, 
    -2.205, -2.17, -2.405, -3.215, -3.525, -3.61, 0.655, 3.6, 5.785, 6.57, 
    6.995, 7.15, 7.53, 7.385, 5.8, 4.335, 4.11, 4.4, 4.24, 4.335, 4.73, 
    4.535, 2.89, 1.555, 0.325, 0.35, 0.845, 0.995, 0.935, 1.355, 1.905, 
    4.155, 4.245, 4.125, 6.345, 5.6, 5.915, 5.98, 5.43, 4.75, 4.135, 3.435, 
    1.83, 1.76, 2.32, 1.64, 0.425, 0.01, -0.145, -0.32, -0.23, -0.18, -0.03, 
    0.285, 0.6, 1.02, 1.555, 2.43, 3, 4.035, 3.705, 3.68, 3.845, 3.64, 2.905, 
    3.01, 3.07, 3.265, 3.21, 2.86, 2.855, 2.865, 2.67, 2.83, 2.345, 1.865, 
    1.64, 1.73, 3.605, 3.61, 3.465, 3.61, 4.065, 4.53, 5.265, 5.195, 5.21, 
    4.105, 3.33, 3.12, 2.525, 1.895, 0.15, 1.09, 0, -0.015, -0.63, 0.365, 
    0.835, -0.315, -0.39, -0.23, 4.315, 6.37, 6.895, 7.54, 8.86, 9.645, 
    9.965, 10.18, 9.68, 7.155, 4.065, 3.22, 3.015, 2.745, 2.37, 2.38, 2.035, 
    2.295, 1.67, 3.37, 4.295, 3.935, 3.145, 3.32, 8.21, 11.115, 11.675, 
    12.655, 13.19, 13.435, 13.86, 13.49, 12.665, 10.17, 7.065, 5.96, 5.635, 
    5.365, 5.86, 5.51, 6.28, 7.3, 6.65, 6.65, 6.48, 6.695, 5.76, 5.82, 10.15, 
    11.875, 13.14, 14.395, 14.8, 14.755, 14.34, 14.805, 13.355, 10.935, 
    8.645, 7.925, 8.335, 8.8, 9.5, 9.395, 9.405, 9.295, 9.275, 8.95, 8.11, 
    6.99, 5.58, 2.68, 3.73, 6.09, 8.08, 7.55, 8.205, 8.445, 7.735, 7.105, 
    3.555, 1.365, 1.605, 0.555, -0.095, -0.245, -0.26, -0.435, -0.365, 
    -0.355, -0.08, -0.255, -0.205, -0.09, -0.065, -0.125, -0.135, 0.01, 
    1.385, 1.325, 2.04, 1.44, 0.56, 1.59, 2, 0.745, -0.065, -1.02, -1.85, 
    -2.13, -2.685, -2.695, -2.875, -2.955, -3.25, -3.665, -3.755, -3.6, 
    -3.76, -3.7, -0.905, -0.065, 1.235, 1.45, 1.37, 1.02, 2.045, 3.05, 2.44, 
    0.715, 0.185, -0.005, -0.605, -0.89, -0.365, -0.47, -0.855, -0.65, 
    -0.475, -0.29, -0.12, -0.145, -1.565, -1.24, -0.695, 0.885, 3.405, 3.905, 
    4.145, 5.08, 5.135, 4.29, 3.015, 1.875, 1.085, 0.55, 0.14, -0.35, -0.775, 
    -1.04, -1.3, -1.82, -2.17, -1.585, -2.265, -1.475, -1.1, -0.55, -0.065, 
    0.42, 1.105, 1.775, 1.865, 1.84, 1.32, 1.39, 1.325, 1.255, 0.875, 1.505, 
    1.655, 0.38, -0.1, -0.275, -0.385, -0.22, 0.45, 0.43, 0.49, 0.57, 0.58, 
    0.53, 0.44, 0.31, 0.385, 0.665, 1.135, 0.99, 1.275, 0.67, 0.04, -1.21, 
    -2.36, -3.435, -3.77, -4.13, -4.62, -4.36, -5.16, -5.175, -5.795, -6.895, 
    -7.15, -7.68, -8.83, -8.525, -5.37, -3.675, -2.575, -2.4, -1.495, -1.24, 
    -1.025, -0.9, -1.645, -3.29, -4.665, -5.31, -6.23, -6.83, -6.85, -6.555, 
    -6.935, -6.27, -5.78, -4.76, -4.385, -5.055, -4.825, -4.195, -2.995, 
    -0.53, 0.425, 0.46, 1.77, 2.12, 1.37, 1.625, 0.675, -0.295, -0.265, 0.47, 
    0.575, 0.845, 1.185, 2.2, 1.26, -1.705, -3.45, -4.61, -5.7, -7.2, -7.61, 
    -7.88, -8.115, -8.325, -8.22, -6.61, -5.275, -5.45, -5.67, -7.43, -8.115, 
    -9.05, -9.905, -9.425, -9.425, -9.975, -10.41, -10.37, -10.525, -10.585, 
    -10.59, -10.185, -10.37, -10.9, -10.375, -10.3, -9.47, -7.345, -4.955, 
    -4.905, -4.81, -3.835, -3.385, -4.11, -4.87, -6.115, -6.84, -7.425, 
    -7.925, -8.435, -8.58, -8.355, -8.895, -9.32, -10.21, -11.555, -10.74, 
    -9.74, -11.12, -11.795, -8.96, -8.105, -6.325, -5.97, -5.05, -4.475, 
    -5.55, -6.345, -7.165, -8.095, -8.82, -9.12, -9.48, -9.46, -9.425, 
    -9.385, -9.26, -8.82, -8.485, -8.135, -7.27, -6.12, -5.78, -4.615, 
    -3.995, -4.02, -4.47, -3.84, -3.655, -3.445, -2.9, -2.355, -2.185, 
    -2.095, -1.985, -1.8, -1.595, -1.53, -1.515, -1.49, -1.565, -1.435, 
    -1.435, -1.68, -1.955, -2.365, -2.435, -2.37, -1.365, -0.055, 0.575, 1.5, 
    3.035, 3.68, 4.335, 4.95, 3.63, 1.775, 0.865, 0.36, 0.275, 0.995, 1.82, 
    1.785, 1.4, 1.36, 1.285, 1.6, 1.835, 1.875, 1.515, 1.73, 3.245, 4.875, 
    5.565, 6.04, 5.82, 5.32, 5.02, 4.055, 4.01, 3.235, 2.145, 1.935, 1.62, 
    1.66, 1.345, 1.35, 0.745, 0.8, 0.725, 0.695, 0.09, 0.1, -0.44, -0.665, 
    1.735, 4.885, 5.61, 6.485, 6.69, 6.055, 6.27, 5.845, 5.125, 3.245, 1.01, 
    0.41, 1.095, 0.325, 0.5, 0.305, 0.655, 1.325, 1.02, 1.255, 0.355, 0.56, 
    0.72, 0.96, 3.15, 5.19, 5.59, 7.01, 7.335, 7.925, 7.875, 7.895, 6.835, 
    4.98, 2.54, 0.655, 0.6, 0.4, 0.27, 0.49, 0.76, 0.82, 1.415, 3.575, 4.175, 
    1.61, 1.81, 1.805, 5.895, 10.93, 11.875, 12.64, 13.65, 14.125, 14.33, 
    13.455, 11.69, 8.375, 6.52, 6.475, 8.25, 8.96, 7.66, 7.7, 7.52, 7.625, 
    7.815, 6.98, 4.965, 3.055, 2.155, 4.905, 7.49, 9.84, 11.135, 12.03, 
    12.36, 11.785, 12.515, 10.92, 10.01, 8.255, 7.295, 6.835, 7.165, 7.89, 
    8.21, 7.47, 6.67, 6.075, 6.055, 5.65, 5.05, 4.79, 4.53, 4.405, 4.635, 
    6.24, 6.61, 6.805, 7.015, 6.83, 6.02, 4.875, 4.105, 3.2, 2.305, 2.36, 
    2.155, 1.6, 1.145, 0.875, 0.415, -0.01, -0.35, -0.21, -0.37, -0.445, 
    -0.4, -0.04, 0.475, 2.315, 3.425, 4.885, 5.01, 3.305, 2.65, 1.91, 2.11, 
    1.01, -0.785, -2.23, -2.46, -2.97, -3.2, -2.71, -2.51, -2.93, -3.775, 
    -4.095, -4.535, -4.84, -6.07, -6.715, -3.515, -0.39, -0.05, -0.225, 0.32, 
    0.97, 1.155, 0.89, 0.04, -2.045, -3.91, -4.535, -4.6, -5.05, -5.16, 
    -4.72, -4.505, -5.255, -6.435, -6.42, -5.605, -5.01, -5.03, -4.77, 
    -2.195, 2.48, 4.08, 5.16, 5.565, 5.865, 6.11, 5.7, 4.06, 1.125, 0.435, 
    1.28, 0.965, 0.3, 1.215, 0.53, 0.51, 1.36, 0.055, -0.23, -0.62, 0, 0.895, 
    0.905, 1.045, 2.225, 3.185, 4.6, 4.88, 5.415, 4.655, 4.425, 3.8, 1.905, 
    -0.445, -1.38, -1.93, -1.92, 0.985, 2.22, 2.435, 1.735, 1.81, 2.32, 
    2.415, 1.915, 0.91, 2.285, 2.85, 5.575, 7.23, 8.69, 8.46, 7.6, 6.61, 6.31, 
    6.02, 5.235, 4.925, 4.94, 4.37, 3.765, 5.105, 5.15, 4.895, 4.455, 3.955, 
    3.905, 3.905, 3.665, 3.23, 2.34, 2.375, 2.05, 0.97, 0.635, -1.855, -2.95, 
    -3.085, -3.63, -4.23, -5.015, -5.825, -6.425, -7.33, -8.405, -8.91, 
    -8.615, -9.645, -10.04, -10.88, -11.45, -11.965, -12.235, -12.515, 
    -12.415, -10.93, -8.25, -6.695, -6.955, -5.96, -7.365, -6.795, -7.075, 
    -7.945, -9.305, -11.035, -11.44, -11.825, -11.58, -12.035, -12.755, 
    -12.61, -11.075, -10.5, -10.245, -9.655, -9.535, -9.825, -9.65, -9.095, 
    -8.31, -7.095, -7.035, -6.855, -7.495, -8.515, -9.36, -9.965, -10.825, 
    -11.33, -11.56, -11.925, -12.32, -12.825, -12.88, -13.815, -14.32, 
    -14.955, -14.53, -14.415, -14.87, -14.375, -14.77, -14.145, -10.085, 
    -9.09, -8.33, -6.735, -7.955, -7.56, -8.015, -9.275, -10.56, -12.09, 
    -12.675, -13.005, -12.425, -11.535, -10.825, -10.895, -10.755, -10.785, 
    -10.695, -10.23, -10.43, -10.04, -9.725, -7.485, -1.285, -0.29, -0.16, 
    -0.38, -0.045, -0.255, 0.37, -1.49, -2.965, -3.435, -3.87, -3.155, 
    -2.305, -2.33, -2.59, -2.8, -1.925, -1.735, -1.4, -2.195, -2.29, -0.96, 
    -2.005, 0.03, 5.11, 6.15, 6.175, 7.57, 7.14, 7.885, 6.83, 4.14, 0.645, 
    -0.96, -0.375, -0.04, -0.23, -0.145, -0.28, -1.02, 0.615, 0.77, 0.62, 
    0.16, 0.315, -0.91, -2.27, -0.615, 4.14, 4.54, 3.83, 3.195, 3.43, 3.36, 
    2.745, 0.845, -0.315, -1.91, -2.33, -2.745, -3.535, -4.07, -5.01, -5.47, 
    -5.905, -7.04, -7.385, -7.685, -7.2, -6.375, -6.535, -5.69, -3.28, 
    -0.525, 0.79, 0.905, 1.02, 1.56, 1.49, -0.495, -2.175, -2.895, -3.095, 
    -3.4, -2.645, -1.965, -2.055, -2.165, -2.97, -4.335, -3.815, -2.18, 0.21, 
    0.665, 0.43, 0.655, 3.58, 3.495, 4.245, 4.465, 4.85, 4.59, 4.26, 3.67, 
    2.045, 1.785, 2.055, 2.625, 2.445, 2.395, 2.105, 1.475, 0.92, -0.795, 
    -2.14, -3.39, -5.35, -5.66, -5.84, -6.37, -6.355, -6.04, -6.16, -6.745, 
    -6.245, -6.955, -7.37, -8, -8.72, -9.125, -9.62, -10.505, -11.24, -11.81, 
    -12.43, -12.6, -13.06, -13.38, -11.865, -10.825, -10.53, -11.27, -10.905, 
    -9.55, -7.595, -4.085, -3.155, -4.43, -5.375, -6.38, -6.51, -6.2, -7.65, 
    -8.285, -8.77, -9.165, -9.735, -10.02, -10.195, -10.51, -10.71, -10.93, 
    -11.065, -11, -11.06, -11.17, -11.32, -11.375, -10.61, -9.92, -8.895, 
    -8.965, -8.75, -8.755, -9.17, -10.595, -10.675, -10.62, -11.175, -11.345, 
    -11.39, -11.695, -11.66, -11.335, -11.495, -12.24, -12.115, -12.18, 
    -12.14, -11.995, -11.935, -10.885, -7.475, -4.39, -2.31, -2.73, -2.565, 
    -1.045, -1.31, -3.53, -4.64, -4.62, -4.335, -5.515, -5.86, -5.425, 
    -5.865, -5.865, -5.38, -5.42, -5.465, -5.11, -4.655, -5, -5.305, -3.68, 
    0.3, 1.87, 2.7, 3.505, 3.69, 4.08, 3.49, 1.735, -0.97, -2.08, -2.675, 
    -3.06, -3.27, -3.89, -3.07, -1.875, -2.305, -2.15, -2.1, -2.715, -2.985, 
    -0.955, -0.215, 0.515, 5.195, 8.785, 9.225, 8.35, 8.725, 7.705, 6.05, 
    3.71, 0.975, -1.16, -2.095, -1.58, -1.835, -0.91, -0.03, -1.605, -1.17, 
    -1.895, -1.175, -1.545, -2.025, -3.73, -3.86, -3.345, 2.315, 3.785, 
    5.015, 4.19, 3.585, 3.145, 2.52, 1.955, -1.575, -3.39, -3.575, -3.205, 
    -2.665, -2.745, -2.525, -2.835, -2.58, -2.665, -2.57, -3.01, -3.335, 
    -3.565, -3.855, -3.535, -2.955, -1.765, 0.75, 1.5, 1.08, 0.455, 0.315, 
    -1.165, -2.665, -3.43, -4.005, -4.715, -5.455, -5.78, -6.79, -7.465, 
    -7.335, -7.735, -7.89, -6.925, -6.36, -5.835, -6.605, -6.105, -2.23, 
    -0.71, 0.665, 1.175, 1.4, 1.33, 0.61, -1.795, -3.185, -4.505, -5.175, 
    -5.71, -6.015, -5.5, -5.5, -5.585, -5.24, -4.56, -4.76, -4.69, -4.35, 
    -4.465, -4.26, -3.565, 1.83, 3.505, 2.76, 2.385, 2.26, 2.495, 1.51, 
    0.325, -1.195, -1.64, -2.145, -2.565, -3.025, -3.54, -3.24, -3.705, 
    -4.01, -4.6, -4.815, -4.81, -4.86, -5.15, -5.755, -5.32, -3.705, -2.425, 
    -1.77, -2.05, -3.41, -4.075, -4.72, -5.075, -5.605, -6.04, -6.7, -7.5, 
    -7.795, -8.12, -8.675, -10.235, -11.22, -11.485, -12.015, -12.63, -13.78, 
    -15.085, -15.58, -14.845, -11.125, -8.695, -6.685, -6.2, -6.495, -6.385, 
    -7.42, -9.66, -11.865, -13.28, -14.14, -14.65, -15.61, -16.54, -16.78, 
    -17.69, -17.96, -18.28, -18.675, -19.345, -19.56, -19.125, -19.805, 
    -19.305, -14.49, -11.81, -11.34, -11.38, -10.775, -10.575, -10.95, 
    -12.405, -14.26, -15.32, -16.83, -15.885, -16.525, -16.755, -16.51, 
    -15.7, -15.335, -15.35, -15.14, -14.785, -14.17, -13.585, -13.835, 
    -14.24, -12.725, -10.805, -9.535, -7.9, -7.18, -6.33, -7.795, -9.215, 
    -10.115, -9.975, -9.47, -9.36, -9.225, -8.995, -9.485, -9.485, -9.63, 
    -10.185, -11.245, -9.905, -9.77, -10.84, -12.165, -12.645, -12.71, 
    -12.485, -11.98, -10.905, -10.755, -11.565, -12.84, -14.165, -15.435, 
    -15.755, -15.655, -16.355, -17.17, -16.77, -16.02, -15.865, -16.38, 
    -17.825, -18.595, -19.02, -19.315, -19.555, -19.755, -19.985, -19.705, 
    -19.19, -18.81, -18.725, -18.26, -18.495, -18.97, -19.66, -20.705, 
    -21.335, -21.745, -22.295, -23.25, -24.245, -24.665, -24.505, -24.485, 
    -24.37, -24.205, -23.345, -22.25, -22.24, -22.17, -22.07, -21.72, 
    -18.895, -19.35, -17.555, -14.885, -12.675, -15.025, -18.625, -17.785, 
    -16.245, -17.095, -16.09, -16.875, -17.51, -18.045, -18.28, -18.3, 
    -18.415, -17.535, -16.975, -17.025, -17.1, -17.755, -18.285, -18.105, 
    -18.125, -17.525, -17.12, -17.48, -18.1, -18.54, -19.775, -20.585, 
    -21.17, -21.385, -21.095, -21.08, -21.235, -20.99, -20.805, -20.515, 
    -20.42, -20.185, -20.075, -20.405, -20.71, -21.015, -20.97, -20.575, 
    -20.225, -19.76, -19.475, -19.22, -19.465, -19.27, -19.115, -19.405, 
    -19.44, -19.37, -19.37, -19.395, -19.415, -19.415, -19.275, -19.17, 
    -19.21, -19.08, -18.99, -18.95, -18.815, -19.28, -18.905, -15.135, 
    -12.275, -11.595, -10.325, -10.455, -11.855, -12.435, -14.485, -15.87, 
    -17.055, -16.975, -16.375, -16.115, -16.07, -16, -15.48, -15.11, -14.535, 
    -14.875, -14.745, -14.215, -13.755, -13.425, -12.825, -10.51, -7.39, 
    -5.575, -4.445, -4.69, -4.975, -6.65, -7.895, -9.725, -11.065, -10.655, 
    -11.37, -10.1, -9.975, -9.885, -9.42, -9.41, -8.945, -8.61, -8.47, 
    -8.175, -7.835, -7.43, -7.385, -7.315, -6.92, -6.52, -6.23, -5.77, -5.79, 
    -6.225, -6.285, -6.125, -5.98, -5.755, -5.645, -5.51, -5.42, -5.425, 
    -5.535, -5.615, -5.5, -5.315, -5.195, -5.08, -5.12, -5.225, -5.365, 
    -5.59, -5.365, -5.44, -5.41, -5.505, -5.91, -6.135, -6.27, -6.38, -6.515, 
    -6.58, -6.55, -6.56, -6.645, -6.965, -7.265, -7.38, -7.825, -7.89, -7.78, 
    -7.7, -7.755, -7.95, -8.075, -8.12, -8.325, -8.255, -7.81, -8.43, -8.73, 
    -8.65, -9.255, -9.505, -9.465, -9.515, -9.92, -10.06, -10.07, -10.025, 
    -9.935, -9.81, -9.62, -8.785, -8.325, -8.485, -8.735, -8.785, -8.92, 
    -5.815, -4.445, -2.155, -2.13, -4.205, -4.08, -5.545, -6.225, -6.72, 
    -6.51, -6.09, -5.84, -5.775, -5.79, -5.185, -5.145, -4.935, -4.48, -4.06, 
    -3.765, -3.84, -4.545, -4.635, -3.765, -2.795, -2.095, -2.21, -2.855, 
    -3.545, -3.3, -3.06, -2.925, -3.525, -3.695, -3.95, -3.685, -3.495, 
    -3.18, -2.925, -3.41, -3.555, -3.325, -3.215, -3.42, -3.67, -3.945, 
    -4.09, -4.305, -4.125, -3.16, -3.65, -3.36, -2.73, -2.61, -3.21, -4.645, 
    -5.35, -5.675, -5.55, -5.51, -5.575, -5.635, -6.055, -6.94, -7.69, 
    -8.405, -9.185, -8.205, -7.705, -7.895, -7.725, -7.58, -6.49, -3.005, 
    -4.335, -3.93, -4.2, -3.965, -5.115, -6.095, -7.21, -7.88, -8.145, 
    -8.285, -8.885, -8.875, -8.96, -9.115, -8.93, -9.305, -9.47, -9.33, 
    -7.835, -7.315, -7.565, -7.18, -6.55, -5.3, -4.76, -4.48, -4.66, -4.61, 
    -4.58, -4.835, -5.255, -5.445, -5.325, -5.35, -5.245, -5.005, -4.79, 
    -4.74, -4.655, -4.06, -3.845, -3.125, -3.29, -2.995, -3.185, -3.31, 
    -2.025, 1.175, 2.505, 3.175, 3.145, 2.57, 1.095, -1.35, -2.875, -3.63, 
    -4.415, -5.305, -5.74, -4.94, -4.63, -4.425, -4.875, -5.035, -4.79, 
    -5.865, -5.805, -5.955, -5.34, -5.38, -2.91, -0.385, -0.27, 0.215, -0.42, 
    -0.215, -1.255, -2.87, -4.465, -5.465, -7.125, -7.495, -6.945, -5.57, 
    -5.24, -4.35, -4.25, -4.575, -4.62, -4.525, -4.58, -5.09, -5.075, -5.31, 
    -5.065, -4.22, -4.815, -5.265, -5.525, -6.25, -6.02, -6.115, -6.55, 
    -6.92, -6.215, -5.89, -5.82, -5.755, -5.795, -6.735, -8.43, -9.43, -8.76, 
    -8.13, -7.59, -7.745, -8.195, -8.035, -7.89, -7.93, -8.515, -8.45, -8.89, 
    -9.35, -10.29, -11.62, -12.92, -13.94, -14.675, -15.21, -16, -16.61, 
    -16.38, -17.19, -17.32, -17.855, -17.57, -18.915, -18.505, -17.815, 
    -18.93, -19.07, -15.53, -13.015, -12.67, -12.56, -12.655, -11.455, 
    -12.965, -14.29, -15.45, -15.815, -15.785, -15.355, -14.63, -14.145, 
    -14.09, -14.285, -14.1, -13.745, -13.875, -14.36, -14.435, -13.25, -12.4, 
    -12.58, -11.29, -8.965, -8.625, -8.975, -9.55, -10.125, -11.08, -11.315, 
    -12.695, -13.315, -13.875, -13.795, -14.37, -14.84, -13.87, -13.465, 
    -13.915, -14.755, -15.205, -15.305, -15.57, -15.355, -15.43, -14.65, 
    -9.12, -4.545, -3, -5.655, -6.365, -6.82, -6.97, -8.125, -10.44, -12.505, 
    -12.785, -12.57, -11.98, -11.945, -12.24, -11.8, -11.285, -10.035, 
    -10.09, -9.615, -10.11, -10.335, -9.92, -10.165, -7.91, -5.725, -5.41, 
    -5.31, -5.18, -5.97, -6.53, -7.595, -8.935, -9.815, -10.375, -10.545, 
    -11.495, -11.895, -12.705, -12.995, -12.85, -13.365, -12.865, -13.145, 
    -13.335, -13.625, -11.99, -12.155, -7.805, -2.85, -2.62, -2.51, -2.495, 
    -2.89, -3.86, -5.75, -8.58, -10.49, -9.89, -9.2, -9.57, -9.025, -9.41, 
    -9.21, -10.37, -10.85, -10.56, -9.405, -9.39, -10.125, -10.545, -9.535, 
    -8.555, -7.765, -8.935, -8.975, -8.225, -8.225, -8.305, -9.36, -10.3, 
    -10.46, -10.32, -10.325, -10.44, -10.57, -10.73, -10.81, -10.83, -10.85, 
    -10.68, -10.515, -10.485, -10.46, -10.375, -10.2, -9.87, -9.71, -9.97, 
    -10.115, -10.29, -10.265, -10.525, -10.655, -10.83, -11.13, -11.32, 
    -11.45, -11.365, -11.41, -11.175, -11, -11.05, -11.16, -11.21, -11.25, 
    -11.325, -11.46, -11.74, -11.78, -11.23, -10.245, -9.775, -9.115, -8.925, 
    -10.265, -10.64, -11.025, -11.22, -11.205, -11.165, -11, -10.64, -10.21, 
    -9.67, -8.725, -7.44, -7.26, -7.165, -6.45, -6.07, -5.98, -5.965, -5.635, 
    -4.63, -3.835, -3.85, -3.82, -4.06, -3.585, -4.02, -4.765, -5.095, -5.26, 
    -5.36, -5, -4.545, -4.355, -4.075, -4.35, -4.48, -4.435, -4.39, -4.57, 
    -4.73, -5.175, -5.51, -6.235, -6.595, -6.35, -6.12, -6.375, -5.735, 
    -6.26, -6.19, -6.82, -7.175, -7.385, -7.775, -8.295, -8.16, -8.425, 
    -8.16, -7.82, -7.76, -7.835, -7.975, -8.065, -8.135, -8.09, -7.875, 
    -7.91, -7.56, -6.925, -5.675, -5.265, -4.71, -4.275, -5.165, -7.075, 
    -7.53, -8.385, -10.07, -11.04, -9.97, -9.465, -9.525, -9.72, -9.175, 
    -8.805, -9.18, -8.68, -9.065, -9.46, -9.745, -8.465, -6.73, -3.945, 
    -0.485, -0.495, -0.645, -2.17, -4.61, -5.76, -6.04, -6.25, -6.28, -5.96, 
    -6.185, -5.615, -5.485, -5.62, -5.33, -5.25, -5.07, -4.695, -4.665, 
    -4.62, -4.345, -4.385, -4.2, -4.09, -4.535, -3.27, -3.08, -3.26, -3.99, 
    -4.615, -5.075, -5.045, -4.375, -4.35, -4.355, -4.49, -4.785, -4.645, 
    -4.725, -4.53, -4.265, -4.075, -3.99, -3.95, -3.695, -3.64, -3.775, 
    -3.84, -3.81, -3.76, -3.865, -4.39, -4.74, -5.52, -6.44, -7.42, -7.99, 
    -8.725, -10.68, -12.035, -12.77, -12.49, -13.635, -15.155, -15.77, 
    -16.06, -16.15, -15.66, -15.92, -15.74, -12.88, -9.905, -6.055, -4.78, 
    -5.285, -5.765, -7.07, -8.32, -10.375, -12.445, -12.86, -12.95, -13.015, 
    -12.6, -12.31, -11.595, -11.38, -11.495, -11.11, -11.01, -10.505, -10.46, 
    -10.64, -10.375, -7.355, -3.06, -0.025, 0.585, -1.085, -1.615, -2.14, 
    -2.935, -4.09, -4.345, -5.01, -4.615, -4.715, -4.73, -4.525, -4.585, 
    -4.71, -5.085, -4.83, -4.06, -4.135, -4.375, -4.645, -5.415, -4.645, 
    -2.545, -1.125, -0.895, -0.94, -1.635, -2.395, -2.705, -3.54, -4.98, 
    -4.475, -4.38, -4.09, -5.535, -5.845, -5.85, -4.81, -4.02, -4.13, -4.63, 
    -5.645, -5.195, -5.64, -5.865, -2.765, 0.66, 1.53, 1.22, 1.9, 1.68, 1.07, 
    -0.37, -1.655, -3.4, -4.36, -4.665, -4.765, -4.8, -4.94, -5.55, -5.315, 
    -5.13, -4.915, -5.165, -5.695, -5.65, -5.645, -5.63, -1.34, 2.43, 3.78, 
    4.19, 3.38, 3.8, 3.395, 1.47, 0.345, -0.085, -0.675, -0.12, -2.305, 
    -4.25, -4.78, -4.225, -4.34, -5.215, -5.575, -2.12, -3.445, -1.35, 
    -0.435, -0.095, 1.43, 1.76, 2.09, 2.54, 2.19, 1.905, 1.185, 1.175, 
    -0.655, -1.435, -2.045, -1.88, -3.135, -3.9, -3.785, -2.76, -2.755, 
    -2.575, -3.11, -4.3, -5.945, -6.455, -6.14, -5.77, -3.155, 0.405, 2.715, 
    2.23, 2.61, 0.42, 1.26, -0.115, -1.685, -2.155, -2.805, -3.24, -3.125, 
    -3.45, -4.3, -4.965, -5.03, -5.665, -5.7, -5.585, -5.795, -5.925, -6.055, 
    -6.155, -5.78, -5.09, -5.12, -4.5, -4.32, -4.195, -4.57, -5.32, -6.03, 
    -6.63, -7.41, -8.055, -8.335, -8.65, -8.58, -8.6, -9.29, -10.37, -10.12, 
    -9.49, -8.435, -8.325, -9.545, -7.535, -6.17, -4.84, -3.28, -2.545, 
    -2.07, -1.18, -1.835, -2.55, -2.56, -2.47, -2.72, -2.68, -3.175, -3.03, 
    -2.35, -2.535, -3.365, -3.07, -3.2, -3.105, -4.345, -3.715, -3.79, 
    -3.585, -1.015, 0.52, 2.87, 3.41, 2.845, 1.565, 1.67, 0.03, -2.025, 
    -2.87, -3.785, -3.61, -3.735, -3.275, -2.905, -3.425, -2.73, -3.705, 
    -3.81, -4.375, -5.085, -6.665, -5.465, -4.25, -1.75, 1.065, 0.805, 1.4, 
    2.235, 2.115, 1.685, -0.19, -2.595, -4.095, -4.015, -3.665, -3.205, 
    -3.03, -2.985, -3.485, -4.155, -4.565, -5.53, -5.695, -4.95, -5.59, 
    -5.92, -5.84, -5.445, -4.705, -4.615, -3.24, -3.86, -3.725, -4.13, -4.04, 
    -4.295, -4.435, -4.19, -4.33, -4.815, -5.005, -5.065, -4.825, -4.8, 
    -4.64, -4.24, -4.485, -4.825, -4.995, -5.245, -5.265, -5.22, -5.775, 
    -5.79, -5.325, -4.55, -5.65, -5.77, -5.91, -7.145, -7.855, -9.365, -8.31, 
    -7.795, -7.275, -7.145, -7.52, -7.775, -7.36, -7.85, -8.25, -8.15, -8.14, 
    -8.6, -8.595, -7.36, -5.85, -4.705, -5.065, -5.045, -5.975, -5.795, 
    -5.55, -6.68, -7.605, -8.11, -7.86, -7.685, -7.485, -7.135, -7.315, 
    -7.36, -7.205, -6.965, -6.82, -6.835, -6.99, -6.895, -6.84, -6.525, 
    -6.02, -5.675, -4.24, -4.675, -4.665, -4.695, -5.27, -6.405, -7.235, 
    -7.1, -7.345, -7.725, -7.48, -7.275, -7.79, -7.68, -7.6, -7.385, -6.56, 
    -5.955, -6.11, -6.545, -6.635, -6.515, -6.17, -5.305, -5.655, -6.005, 
    -6.695, -7.035, -7.16, -7.205, -7.37, -7.59, -7.7, -7.82, -8.26, -8.495, 
    -8.565, -8.605, -8.81, -9.19, -9.41, -9.475, -9.51, -9.555, -9.64, -9.5, 
    -9.35, -9.2, -9.22, -9.44, -9.615, -9.78, -9.78, -9.685, -9.65, -9.625, 
    -9.6, -9.625, -9.74, -9.875, -9.965, -10.075, -10.175, -10.23, -10.215, 
    -10.255, -10.31, -10.31, -10.375, -10.22, -9.755, -8.63, -7.215, -8.505, 
    -9.28, -9.46, -10.105, -10.5, -10.91, -11.29, -11.585, -11.655, -11.925, 
    -12.14, -12.165, -11.54, -11.055, -11.17, -11.26, -10.815, -10.49, 
    -10.505, -10.025, -9.39, -9.115, -8.83, -8.345, -6.725, -6.045, -5.165, 
    -5.88, -7.2, -7.63, -7.795, -8.485, -10.6, -11.19, -9.17, -8.75, -9.605, 
    -10.255, -10.735, -10.06, -8.325, -6.455, -6.355, -6.43, -5.34, -3.955, 
    -2.875, -3.755, -3.085, -2.67, -2.3, -3.165, -4.445, -5.105, -5.345, 
    -5.525, -6.06, -6.5, -7.16, -7.35, -7.11, -8.16, -8.68, -8.495, -8.6, 
    -8.165, -7.945, -8.435, -6.715, -4.175, -2.98, -2.245, -2.635, -2.99, 
    -3.59, -4.015, -5.26, -6.64, -6.955, -6.945, -6.925, -6.8, -7.245, -7.65, 
    -8, -8.105, -8.07, -7.99, -8.055, -8.935, -9.44, -9.425, -6.345, -4.485, 
    -3.795, -3.12, -2.88, -2.25, -2.125, -3.3, -5.79, -7.66, -8.255, -8.985, 
    -9.48, -9.625, -10.43, -10.325, -9.5, -10.63, -10.7, -10.325, -10.52, 
    -10.815, -10.675, -10.165, -6.18, -3.14, -1.37, -1.145, -0.9, -0.62, 
    -0.66, -3.105, -4.88, -6.73, -6.945, -7.765, -8.805, -8.975, -8.825, 
    -8.2, -7.88, -9.39, -8.385, -8.9, -7.305, -7.37, -9.75, -9.985, -6.56, 
    -1.025, 1.22, 1.44, 0.785, 0.615, 0.5, -1.65, -3.605, -4.805, -5.71, 
    -5.435, -5.24, -5.53, -5.61, -5.725, -6.06, -6.46, -6.985, -7.275, 
    -7.265, -7.285, -7.25, -7.255, -7.085, -6.685, -6.695, -6.635, -6.77, 
    -6.92, -6.815, -7.225, -7.32, -7.365, -7.32, -7.345, -7.475, -7.72, 
    -7.725, -7.9, -8.01, -8.005, -8.005, -8.155, -8.295, -8.405, -8.615, 
    -8.675, -8.375, -7.33, -6.57, -6.145, -7.515, -6.66, -5.42, -6.335, 
    -7.645, -8.825, -9.915, -11.955, -11.91, -11.31, -10.255, -10.925, 
    -10.965, -10.295, -9.375, -9.245, -9.375, -9.755, -10.95, -10.68, -6.425, 
    -0.755, -0.125, -1.15, -2.785, -3.34, -3.385, -3.89, -4.725, -6.705, 
    -7.995, -7.465, -7.3, -7.64, -9.24, -9.84, -10.31, -9.99, -9.83, -9.6, 
    -9.3, -8.495, -7.625, -6.185, -4.885, -5.4, -4.21, -1.24, -1.065, -1.255, 
    -1.425, -2.215, -3.815, -5.24, -5.98, -5.975, -6.325, -6.35, -6.46, 
    -6.48, -6.93, -7.535, -7.795, -8.035, -8.045, -7.93, -8.735, -8.93, 
    -7.295, -6.155, -6.31, -5.095, -4.445, -5.165, -6.095, -5.32, -6.735, 
    -8.38, -9.31, -9.57, -9.25, -9.895, -9.365, -8.545, -8.21, -7.295, -6.67, 
    -7.195, -6.61, -6.67, -6.725, -6.145, -5.555, -5.355, -4.36, -3.695, 
    -4.14, -4.485, -4.5, -4.57, -4.555, -4.615, -4.52, -4.37, -4.4, -4.33, 
    -4.315, -4.195, -4.16, -4.23, -4.41, -4.47, -4.605, -4.95, -5.225, -4.84, 
    -4, -3.795, -2.98, -1.985, -2.375, -2.63, -2.42, -2.535, -4.08, -6.485, 
    -6.71, -5.935, -6.07, -6.475, -6.465, -6.67, -6.925, -7.095, -7.7, -7.6, 
    -7.435, -7.48, -7.89, -8.11, -8.09, -8, -7.58, -7.225, -6.825, -6.825, 
    -6.71, -6.68, -7.045, -8.085, -8.965, -9.575, -9.685, -9.85, -10.19, 
    -10.47, -11.075, -11.385, -11.22, -12.165, -12.885, -14.19, -14.465, 
    -13.165, -6.15, -5.99, -6.675, -5.78, -4.725, -6.39, -7.43, -8.135, 
    -8.98, -10.35, -10.75, -11.035, -12.695, -13.41, -13.825, -14.255, 
    -14.295, -14.6, -15.105, -13.685, -12.32, -11.06, -11.32, -10.655, -9.62, 
    -9.305, -8.37, -8.195, -6.635, -8.045, -7.84, -7.43, -8.675, -11.25, 
    -13.195, -11.835, -12.225, -12.505, -11.32, -11.215, -10.7, -10.465, 
    -10.26, -9.855, -9.795, -9.725, -9.865, -9.715, -8.72, -8.1, -7.4, -6.72, 
    -6.94, -8.03, -7.95, -7.94, -8.505, -8.735, -8.84, -8.865, -9.165, -9.31, 
    -9.26, -9.06, -9.1, -9.045, -8.615, -8.56, -8.64, -8.805, -8.88, -8.76, 
    -8.4, -7.845, -7.49, -7.125, -7.01, -6.955, -6.95, -6.745, -6.995, -7.18, 
    -7.28, -7.07, -7.095, -7.025, -6.625, -6.395, -6.305, -6.3, -6.215, 
    -6.22, -6.33, -6.355, -6.22, -5.985, -5.475, -5.3, -5.195, -4.985, -4.92, 
    -4.855, -5.115, -5.4, -5.455, -5.76, -5.695, -5.47, -5.305, -5.165, 
    -5.085, -5.23, -5.325, -5.285, -5.295, -5.315, -5.375, -5.275, -5.255, 
    -5.175, -4.885, -4.745, -4.825, -4.745, -4.745, -4.535, -5.295, -5.79, 
    -6.865, -8.16, -8.745, -9.715, -10.79, -9.655, -10.88,
  -7.355, -7.545, -6.75, -6.6, -6.515, -6.545, -7.34, -7.17, -5.715, -3.385, 
    -2.5, -2.31, -2.12, -1.97, -1.89, -2.04, -2.135, -3.33, -4.08, -4.8, 
    -5.035, -5.04, -4.9, -5.815, -5.1, -5.15, -5.315, -5.8, -6.785, -6.35, 
    -5.995, -4.845, -0.33, 1.05, 2.065, 2.82, 3.24, 4.18, 5.065, 4.925, 
    3.445, 2.475, 0.415, -2.325, -2.92, -3.28, -3.53, -2.68, -1.465, -2.74, 
    -1.81, -1.145, -0.18, -0.495, -0.52, 0.235, 1.205, 2.535, 2.73, 3.665, 
    4.295, 4.175, 4.94, 4.9, 4.45, 4.64, 2.975, 2.725, 2.615, 2.685, 2.435, 
    1.81, 0.91, 0.205, -0.235, -0.47, -0.515, -0.64, -0.845, -1.78, -2.05, 
    -1.92, -2.125, -1.23, -1.25, -1.145, -1.6, -1.23, -1.585, -1.585, -2.3, 
    -3.15, -3.33, -3.36, -3.455, -3.855, -4.075, -4.75, -4.96, -5.165, 
    -5.515, -5.835, -6.545, -6.57, -5.72, -5.005, -4.595, -4.815, -3.385, 
    -3.49, -4.83, -4.685, -4.665, -4.815, -4.99, -5.62, -5.855, -6.195, 
    -6.57, -7.72, -6.98, -8.075, -8.33, -7.45, -7.99, -9.205, -9.06, -7.505, 
    -3.675, -0.52, -1.075, 0.005, 0.47, 0.59, 1.325, 1.63, 1.59, -0.02, 
    -1.915, -3.25, -3.25, -2.425, -4.04, -5.65, -5.835, -5.745, -5.095, 
    -5.94, -6.22, -4.83, -5.01, -4.02, 1.03, 3.93, 4.6, 4.285, 5.385, 5.39, 
    5.855, 5.045, 3.88, 2.25, -0.07, -1.25, -1.275, -1.83, -2.23, -2.965, 
    -3.6, -4.115, -3.435, -3.18, -3.76, -4.225, -3.655, -3.03, -2.51, -2.165, 
    0.25, 0.005, 0.1, -0.37, -0.09, 0.575, -0.515, -1.49, -1.795, -1.965, 
    -2.835, -2.945, -2.88, -3.1, -3.305, -3.18, -3.02, -3.015, -2.87, -2.635, 
    -2.615, -2.5, -2.25, -1.475, -1.045, -0.975, -0.885, -0.44, 0.04, 0.575, 
    0.585, 0.22, -0.6, -1.41, -1.905, -2.355, -2.885, -3.295, -3.56, -3.7, 
    -3.8, -4.255, -4.765, -5.17, -5.03, -5.185, -4.64, -3.875, -3.515, 
    -1.445, -0.825, -1.09, -1.695, -2.995, -3.1, -3.2, -3.325, -3.35, -3.39, 
    -3.75, -3.445, -3.285, -3.715, -4.055, -3.645, -3.545, -3.24, -2.81, 
    -2.575, -2.42, -2.11, -1.765, -1.535, -1.51, -1.54, -1.775, -1.7, -0.625, 
    -0.39, -0.87, -1.65, -2.055, -2.42, -2.41, -2.55, -2.84, -2.545, -2.04, 
    -2.205, -2.17, -2.405, -3.215, -3.525, -3.61, 0.655, 3.6, 5.785, 6.57, 
    6.995, 7.15, 7.53, 7.385, 5.8, 4.335, 4.11, 4.4, 4.24, 4.335, 4.73, 
    4.535, 2.89, 1.555, 0.325, 0.35, 0.845, 0.995, 0.935, 1.355, 1.905, 
    4.155, 4.245, 4.125, 6.345, 5.6, 5.915, 5.98, 5.43, 4.75, 4.135, 3.435, 
    1.83, 1.76, 2.32, 1.64, 0.425, 0.01, -0.145, -0.32, -0.23, -0.18, -0.03, 
    0.285, 0.6, 1.02, 1.555, 2.43, 3, 4.035, 3.705, 3.68, 3.845, 3.64, 2.905, 
    3.01, 3.07, 3.265, 3.21, 2.86, 2.855, 2.865, 2.67, 2.83, 2.345, 1.865, 
    1.64, 1.73, 3.605, 3.61, 3.465, 3.61, 4.065, 4.53, 5.265, 5.195, 5.21, 
    4.105, 3.33, 3.12, 2.525, 1.895, 0.15, 1.09, 0, -0.015, -0.63, 0.365, 
    0.835, -0.315, -0.39, -0.23, 4.315, 6.37, 6.895, 7.54, 8.86, 9.645, 
    9.965, 10.18, 9.68, 7.155, 4.065, 3.22, 3.015, 2.745, 2.37, 2.38, 2.035, 
    2.295, 1.67, 3.37, 4.295, 3.935, 3.145, 3.32, 8.21, 11.115, 11.675, 
    12.655, 13.19, 13.435, 13.86, 13.49, 12.665, 10.17, 7.065, 5.96, 5.635, 
    5.365, 5.86, 5.51, 6.28, 7.3, 6.65, 6.65, 6.48, 6.695, 5.76, 5.82, 10.15, 
    11.875, 13.14, 14.395, 14.8, 14.755, 14.34, 14.805, 13.355, 10.935, 
    8.645, 7.925, 8.335, 8.8, 9.5, 9.395, 9.405, 9.295, 9.275, 8.95, 8.11, 
    6.99, 5.58, 2.68, 3.73, 6.09, 8.08, 7.55, 8.205, 8.445, 7.735, 7.105, 
    3.555, 1.365, 1.605, 0.555, -0.095, -0.245, -0.26, -0.435, -0.365, 
    -0.355, -0.08, -0.255, -0.205, -0.09, -0.065, -0.125, -0.135, 0.01, 
    1.385, 1.325, 2.04, 1.44, 0.56, 1.59, 2, 0.745, -0.065, -1.02, -1.85, 
    -2.13, -2.685, -2.695, -2.875, -2.955, -3.25, -3.665, -3.755, -3.6, 
    -3.76, -3.7, -0.905, -0.065, 1.235, 1.45, 1.37, 1.02, 2.045, 3.05, 2.44, 
    0.715, 0.185, -0.005, -0.605, -0.89, -0.365, -0.47, -0.855, -0.65, 
    -0.475, -0.29, -0.12, -0.145, -1.565, -1.24, -0.695, 0.885, 3.405, 3.905, 
    4.145, 5.08, 5.135, 4.29, 3.015, 1.875, 1.085, 0.55, 0.14, -0.35, -0.775, 
    -1.04, -1.3, -1.82, -2.17, -1.585, -2.265, -1.475, -1.1, -0.55, -0.065, 
    0.42, 1.105, 1.775, 1.865, 1.84, 1.32, 1.39, 1.325, 1.255, 0.875, 1.505, 
    1.655, 0.38, -0.1, -0.275, -0.385, -0.22, 0.45, 0.43, 0.49, 0.57, 0.58, 
    0.53, 0.44, 0.31, 0.385, 0.665, 1.135, 0.99, 1.275, 0.67, 0.04, -1.21, 
    -2.36, -3.435, -3.77, -4.13, -4.62, -4.36, -5.16, -5.175, -5.795, -6.895, 
    -7.15, -7.68, -8.83, -8.525, -5.37, -3.675, -2.575, -2.4, -1.495, -1.24, 
    -1.025, -0.9, -1.645, -3.29, -4.665, -5.31, -6.23, -6.83, -6.85, -6.555, 
    -6.935, -6.27, -5.78, -4.76, -4.385, -5.055, -4.825, -4.195, -2.995, 
    -0.53, 0.425, 0.46, 1.77, 2.12, 1.37, 1.625, 0.675, -0.295, -0.265, 0.47, 
    0.575, 0.845, 1.185, 2.2, 1.26, -1.705, -3.45, -4.61, -5.7, -7.2, -7.61, 
    -7.88, -8.115, -8.325, -8.22, -6.61, -5.275, -5.45, -5.67, -7.43, -8.115, 
    -9.05, -9.905, -9.425, -9.425, -9.975, -10.41, -10.37, -10.525, -10.585, 
    -10.59, -10.185, -10.37, -10.9, -10.375, -10.3, -9.47, -7.345, -4.955, 
    -4.905, -4.81, -3.835, -3.385, -4.11, -4.87, -6.115, -6.84, -7.425, 
    -7.925, -8.435, -8.58, -8.355, -8.895, -9.32, -10.21, -11.555, -10.74, 
    -9.74, -11.12, -11.795, -8.96, -8.105, -6.325, -5.97, -5.05, -4.475, 
    -5.55, -6.345, -7.165, -8.095, -8.82, -9.12, -9.48, -9.46, -9.425, 
    -9.385, -9.26, -8.82, -8.485, -8.135, -7.27, -6.12, -5.78, -4.615, 
    -3.995, -4.02, -4.47, -3.84, -3.655, -3.445, -2.9, -2.355, -2.185, 
    -2.095, -1.985, -1.8, -1.595, -1.53, -1.515, -1.49, -1.565, -1.435, 
    -1.435, -1.68, -1.955, -2.365, -2.435, -2.37, -1.365, -0.055, 0.575, 1.5, 
    3.035, 3.68, 4.335, 4.95, 3.63, 1.775, 0.865, 0.36, 0.275, 0.995, 1.82, 
    1.785, 1.4, 1.36, 1.285, 1.6, 1.835, 1.875, 1.515, 1.73, 3.245, 4.875, 
    5.565, 6.04, 5.82, 5.32, 5.02, 4.055, 4.01, 3.235, 2.145, 1.935, 1.62, 
    1.66, 1.345, 1.35, 0.745, 0.8, 0.725, 0.695, 0.09, 0.1, -0.44, -0.665, 
    1.735, 4.885, 5.61, 6.485, 6.69, 6.055, 6.27, 5.845, 5.125, 3.245, 1.01, 
    0.41, 1.095, 0.325, 0.5, 0.305, 0.655, 1.325, 1.02, 1.255, 0.355, 0.56, 
    0.72, 0.96, 3.15, 5.19, 5.59, 7.01, 7.335, 7.925, 7.875, 7.895, 6.835, 
    4.98, 2.54, 0.655, 0.6, 0.4, 0.27, 0.49, 0.76, 0.82, 1.415, 3.575, 4.175, 
    1.61, 1.81, 1.805, 5.895, 10.93, 11.875, 12.64, 13.65, 14.125, 14.33, 
    13.455, 11.69, 8.375, 6.52, 6.475, 8.25, 8.96, 7.66, 7.7, 7.52, 7.625, 
    7.815, 6.98, 4.965, 3.055, 2.155, 4.905, 7.49, 9.84, 11.135, 12.03, 
    12.36, 11.785, 12.515, 10.92, 10.01, 8.255, 7.295, 6.835, 7.165, 7.89, 
    8.21, 7.47, 6.67, 6.075, 6.055, 5.65, 5.05, 4.79, 4.53, 4.405, 4.635, 
    6.24, 6.61, 6.805, 7.015, 6.83, 6.02, 4.875, 4.105, 3.2, 2.305, 2.36, 
    2.155, 1.6, 1.145, 0.875, 0.415, -0.01, -0.35, -0.21, -0.37, -0.445, 
    -0.4, -0.04, 0.475, 2.315, 3.425, 4.885, 5.01, 3.305, 2.65, 1.91, 2.11, 
    1.01, -0.785, -2.23, -2.46, -2.97, -3.2, -2.71, -2.51, -2.93, -3.775, 
    -4.095, -4.535, -4.84, -6.07, -6.715, -3.515, -0.39, -0.05, -0.225, 0.32, 
    0.97, 1.155, 0.89, 0.04, -2.045, -3.91, -4.535, -4.6, -5.05, -5.16, 
    -4.72, -4.505, -5.255, -6.435, -6.42, -5.605, -5.01, -5.03, -4.77, 
    -2.195, 2.48, 4.08, 5.16, 5.565, 5.865, 6.11, 5.7, 4.06, 1.125, 0.435, 
    1.28, 0.965, 0.3, 1.215, 0.53, 0.51, 1.36, 0.055, -0.23, -0.62, 0, 0.895, 
    0.905, 1.045, 2.225, 3.185, 4.6, 4.88, 5.415, 4.655, 4.425, 3.8, 1.905, 
    -0.445, -1.38, -1.93, -1.92, 0.985, 2.22, 2.435, 1.735, 1.81, 2.32, 
    2.415, 1.915, 0.91, 2.285, 2.85, 5.575, 7.23, 8.69, 8.46, 7.6, 6.61, 6.31, 
    6.02, 5.235, 4.925, 4.94, 4.37, 3.765, 5.105, 5.15, 4.895, 4.455, 3.955, 
    3.905, 3.905, 3.665, 3.23, 2.34, 2.375, 2.05, 0.97, 0.635, -1.855, -2.95, 
    -3.085, -3.63, -4.23, -5.015, -5.825, -6.425, -7.33, -8.405, -8.91, 
    -8.615, -9.645, -10.04, -10.88, -11.45, -11.965, -12.235, -12.515, 
    -12.415, -10.93, -8.25, -6.695, -6.955, -5.96, -7.365, -6.795, -7.075, 
    -7.945, -9.305, -11.035, -11.44, -11.825, -11.58, -12.035, -12.755, 
    -12.61, -11.075, -10.5, -10.245, -9.655, -9.535, -9.825, -9.65, -9.095, 
    -8.31, -7.095, -7.035, -6.855, -7.495, -8.515, -9.36, -9.965, -10.825, 
    -11.33, -11.56, -11.925, -12.32, -12.825, -12.88, -13.815, -14.32, 
    -14.955, -14.53, -14.415, -14.87, -14.375, -14.77, -14.145, -10.085, 
    -9.09, -8.33, -6.735, -7.955, -7.56, -8.015, -9.275, -10.56, -12.09, 
    -12.675, -13.005, -12.425, -11.535, -10.825, -10.895, -10.755, -10.785, 
    -10.695, -10.23, -10.43, -10.04, -9.725, -7.485, -1.285, -0.29, -0.16, 
    -0.38, -0.045, -0.255, 0.37, -1.49, -2.965, -3.435, -3.87, -3.155, 
    -2.305, -2.33, -2.59, -2.8, -1.925, -1.735, -1.4, -2.195, -2.29, -0.96, 
    -2.005, 0.03, 5.11, 6.15, 6.175, 7.57, 7.14, 7.885, 6.83, 4.14, 0.645, 
    -0.96, -0.375, -0.04, -0.23, -0.145, -0.28, -1.02, 0.615, 0.77, 0.62, 
    0.16, 0.315, -0.91, -2.27, -0.615, 4.14, 4.54, 3.83, 3.195, 3.43, 3.36, 
    2.745, 0.845, -0.315, -1.91, -2.33, -2.745, -3.535, -4.07, -5.01, -5.47, 
    -5.905, -7.04, -7.385, -7.685, -7.2, -6.375, -6.535, -5.69, -3.28, 
    -0.525, 0.79, 0.905, 1.02, 1.56, 1.49, -0.495, -2.175, -2.895, -3.095, 
    -3.4, -2.645, -1.965, -2.055, -2.165, -2.97, -4.335, -3.815, -2.18, 0.21, 
    0.665, 0.43, 0.655, 3.58, 3.495, 4.245, 4.465, 4.85, 4.59, 4.26, 3.67, 
    2.045, 1.785, 2.055, 2.625, 2.445, 2.395, 2.105, 1.475, 0.92, -0.795, 
    -2.14, -3.39, -5.35, -5.66, -5.84, -6.37, -6.355, -6.04, -6.16, -6.745, 
    -6.245, -6.955, -7.37, -8, -8.72, -9.125, -9.62, -10.505, -11.24, -11.81, 
    -12.43, -12.6, -13.06, -13.38, -11.865, -10.825, -10.53, -11.27, -10.905, 
    -9.55, -7.595, -4.085, -3.155, -4.43, -5.375, -6.38, -6.51, -6.2, -7.65, 
    -8.285, -8.77, -9.165, -9.735, -10.02, -10.195, -10.51, -10.71, -10.93, 
    -11.065, -11, -11.06, -11.17, -11.32, -11.375, -10.61, -9.92, -8.895, 
    -8.965, -8.75, -8.755, -9.17, -10.595, -10.675, -10.62, -11.175, -11.345, 
    -11.39, -11.695, -11.66, -11.335, -11.495, -12.24, -12.115, -12.18, 
    -12.14, -11.995, -11.935, -10.885, -7.475, -4.39, -2.31, -2.73, -2.565, 
    -1.045, -1.31, -3.53, -4.64, -4.62, -4.335, -5.515, -5.86, -5.425, 
    -5.865, -5.865, -5.38, -5.42, -5.465, -5.11, -4.655, -5, -5.305, -3.68, 
    0.3, 1.87, 2.7, 3.505, 3.69, 4.08, 3.49, 1.735, -0.97, -2.08, -2.675, 
    -3.06, -3.27, -3.89, -3.07, -1.875, -2.305, -2.15, -2.1, -2.715, -2.985, 
    -0.955, -0.215, 0.515, 5.195, 8.785, 9.225, 8.35, 8.725, 7.705, 6.05, 
    3.71, 0.975, -1.16, -2.095, -1.58, -1.835, -0.91, -0.03, -1.605, -1.17, 
    -1.895, -1.175, -1.545, -2.025, -3.73, -3.86, -3.345, 2.315, 3.785, 
    5.015, 4.19, 3.585, 3.145, 2.52, 1.955, -1.575, -3.39, -3.575, -3.205, 
    -2.665, -2.745, -2.525, -2.835, -2.58, -2.665, -2.57, -3.01, -3.335, 
    -3.565, -3.855, -3.535, -2.955, -1.765, 0.75, 1.5, 1.08, 0.455, 0.315, 
    -1.165, -2.665, -3.43, -4.005, -4.715, -5.455, -5.78, -6.79, -7.465, 
    -7.335, -7.735, -7.89, -6.925, -6.36, -5.835, -6.605, -6.105, -2.23, 
    -0.71, 0.665, 1.175, 1.4, 1.33, 0.61, -1.795, -3.185, -4.505, -5.175, 
    -5.71, -6.015, -5.5, -5.5, -5.585, -5.24, -4.56, -4.76, -4.69, -4.35, 
    -4.465, -4.26, -3.565, 1.83, 3.505, 2.76, 2.385, 2.26, 2.495, 1.51, 
    0.325, -1.195, -1.64, -2.145, -2.565, -3.025, -3.54, -3.24, -3.705, 
    -4.01, -4.6, -4.815, -4.81, -4.86, -5.15, -5.755, -5.32, -3.705, -2.425, 
    -1.77, -2.05, -3.41, -4.075, -4.72, -5.075, -5.605, -6.04, -6.7, -7.5, 
    -7.795, -8.12, -8.675, -10.235, -11.22, -11.485, -12.015, -12.63, -13.78, 
    -15.085, -15.58, -14.845, -11.125, -8.695, -6.685, -6.2, -6.495, -6.385, 
    -7.42, -9.66, -11.865, -13.28, -14.14, -14.65, -15.61, -16.54, -16.78, 
    -17.69, -17.96, -18.28, -18.675, -19.345, -19.56, -19.125, -19.805, 
    -19.305, -14.49, -11.81, -11.34, -11.38, -10.775, -10.575, -10.95, 
    -12.405, -14.26, -15.32, -16.83, -15.885, -16.525, -16.755, -16.51, 
    -15.7, -15.335, -15.35, -15.14, -14.785, -14.17, -13.585, -13.835, 
    -14.24, -12.725, -10.805, -9.535, -7.9, -7.18, -6.33, -7.795, -9.215, 
    -10.115, -9.975, -9.47, -9.36, -9.225, -8.995, -9.485, -9.485, -9.63, 
    -10.185, -11.245, -9.905, -9.77, -10.84, -12.165, -12.645, -12.71, 
    -12.485, -11.98, -10.905, -10.755, -11.565, -12.84, -14.165, -15.435, 
    -15.755, -15.655, -16.355, -17.17, -16.77, -16.02, -15.865, -16.38, 
    -17.825, -18.595, -19.02, -19.315, -19.555, -19.755, -19.985, -19.705, 
    -19.19, -18.81, -18.725, -18.26, -18.495, -18.97, -19.66, -20.705, 
    -21.335, -21.745, -22.295, -23.25, -24.245, -24.665, -24.505, -24.485, 
    -24.37, -24.205, -23.345, -22.25, -22.24, -22.17, -22.07, -21.72, 
    -18.895, -19.35, -17.555, -14.885, -12.675, -15.025, -18.625, -17.785, 
    -16.245, -17.095, -16.09, -16.875, -17.51, -18.045, -18.28, -18.3, 
    -18.415, -17.535, -16.975, -17.025, -17.1, -17.755, -18.285, -18.105, 
    -18.125, -17.525, -17.12, -17.48, -18.1, -18.54, -19.775, -20.585, 
    -21.17, -21.385, -21.095, -21.08, -21.235, -20.99, -20.805, -20.515, 
    -20.42, -20.185, -20.075, -20.405, -20.71, -21.015, -20.97, -20.575, 
    -20.225, -19.76, -19.475, -19.22, -19.465, -19.27, -19.115, -19.405, 
    -19.44, -19.37, -19.37, -19.395, -19.415, -19.415, -19.275, -19.17, 
    -19.21, -19.08, -18.99, -18.95, -18.815, -19.28, -18.905, -15.135, 
    -12.275, -11.595, -10.325, -10.455, -11.855, -12.435, -14.485, -15.87, 
    -17.055, -16.975, -16.375, -16.115, -16.07, -16, -15.48, -15.11, -14.535, 
    -14.875, -14.745, -14.215, -13.755, -13.425, -12.825, -10.51, -7.39, 
    -5.575, -4.445, -4.69, -4.975, -6.65, -7.895, -9.725, -11.065, -10.655, 
    -11.37, -10.1, -9.975, -9.885, -9.42, -9.41, -8.945, -8.61, -8.47, 
    -8.175, -7.835, -7.43, -7.385, -7.315, -6.92, -6.52, -6.23, -5.77, -5.79, 
    -6.225, -6.285, -6.125, -5.98, -5.755, -5.645, -5.51, -5.42, -5.425, 
    -5.535, -5.615, -5.5, -5.315, -5.195, -5.08, -5.12, -5.225, -5.365, 
    -5.59, -5.365, -5.44, -5.41, -5.505, -5.91, -6.135, -6.27, -6.38, -6.515, 
    -6.58, -6.55, -6.56, -6.645, -6.965, -7.265, -7.38, -7.825, -7.89, -7.78, 
    -7.7, -7.755, -7.95, -8.075, -8.12, -8.325, -8.255, -7.81, -8.43, -8.73, 
    -8.65, -9.255, -9.505, -9.465, -9.515, -9.92, -10.06, -10.07, -10.025, 
    -9.935, -9.81, -9.62, -8.785, -8.325, -8.485, -8.735, -8.785, -8.92, 
    -5.815, -4.445, -2.155, -2.13, -4.205, -4.08, -5.545, -6.225, -6.72, 
    -6.51, -6.09, -5.84, -5.775, -5.79, -5.185, -5.145, -4.935, -4.48, -4.06, 
    -3.765, -3.84, -4.545, -4.635, -3.765, -2.795, -2.095, -2.21, -2.855, 
    -3.545, -3.3, -3.06, -2.925, -3.525, -3.695, -3.95, -3.685, -3.495, 
    -3.18, -2.925, -3.41, -3.555, -3.325, -3.215, -3.42, -3.67, -3.945, 
    -4.09, -4.305, -4.125, -3.16, -3.65, -3.36, -2.73, -2.61, -3.21, -4.645, 
    -5.35, -5.675, -5.55, -5.51, -5.575, -5.635, -6.055, -6.94, -7.69, 
    -8.405, -9.185, -8.205, -7.705, -7.895, -7.725, -7.58, -6.49, -3.005, 
    -4.335, -3.93, -4.2, -3.965, -5.115, -6.095, -7.21, -7.88, -8.145, 
    -8.285, -8.885, -8.875, -8.96, -9.115, -8.93, -9.305, -9.47, -9.33, 
    -7.835, -7.315, -7.565, -7.18, -6.55, -5.3, -4.76, -4.48, -4.66, -4.61, 
    -4.58, -4.835, -5.255, -5.445, -5.325, -5.35, -5.245, -5.005, -4.79, 
    -4.74, -4.655, -4.06, -3.845, -3.125, -3.29, -2.995, -3.185, -3.31, 
    -2.025, 1.175, 2.505, 3.175, 3.145, 2.57, 1.095, -1.35, -2.875, -3.63, 
    -4.415, -5.305, -5.74, -4.94, -4.63, -4.425, -4.875, -5.035, -4.79, 
    -5.865, -5.805, -5.955, -5.34, -5.38, -2.91, -0.385, -0.27, 0.215, -0.42, 
    -0.215, -1.255, -2.87, -4.465, -5.465, -7.125, -7.495, -6.945, -5.57, 
    -5.24, -4.35, -4.25, -4.575, -4.62, -4.525, -4.58, -5.09, -5.075, -5.31, 
    -5.065, -4.22, -4.815, -5.265, -5.525, -6.25, -6.02, -6.115, -6.55, 
    -6.92, -6.215, -5.89, -5.82, -5.755, -5.795, -6.735, -8.43, -9.43, -8.76, 
    -8.13, -7.59, -7.745, -8.195, -8.035, -7.89, -7.93, -8.515, -8.45, -8.89, 
    -9.35, -10.29, -11.62, -12.92, -13.94, -14.675, -15.21, -16, -16.61, 
    -16.38, -17.19, -17.32, -17.855, -17.57, -18.915, -18.505, -17.815, 
    -18.93, -19.07, -15.53, -13.015, -12.67, -12.56, -12.655, -11.455, 
    -12.965, -14.29, -15.45, -15.815, -15.785, -15.355, -14.63, -14.145, 
    -14.09, -14.285, -14.1, -13.745, -13.875, -14.36, -14.435, -13.25, -12.4, 
    -12.58, -11.29, -8.965, -8.625, -8.975, -9.55, -10.125, -11.08, -11.315, 
    -12.695, -13.315, -13.875, -13.795, -14.37, -14.84, -13.87, -13.465, 
    -13.915, -14.755, -15.205, -15.305, -15.57, -15.355, -15.43, -14.65, 
    -9.12, -4.545, -3, -5.655, -6.365, -6.82, -6.97, -8.125, -10.44, -12.505, 
    -12.785, -12.57, -11.98, -11.945, -12.24, -11.8, -11.285, -10.035, 
    -10.09, -9.615, -10.11, -10.335, -9.92, -10.165, -7.91, -5.725, -5.41, 
    -5.31, -5.18, -5.97, -6.53, -7.595, -8.935, -9.815, -10.375, -10.545, 
    -11.495, -11.895, -12.705, -12.995, -12.85, -13.365, -12.865, -13.145, 
    -13.335, -13.625, -11.99, -12.155, -7.805, -2.85, -2.62, -2.51, -2.495, 
    -2.89, -3.86, -5.75, -8.58, -10.49, -9.89, -9.2, -9.57, -9.025, -9.41, 
    -9.21, -10.37, -10.85, -10.56, -9.405, -9.39, -10.125, -10.545, -9.535, 
    -8.555, -7.765, -8.935, -8.975, -8.225, -8.225, -8.305, -9.36, -10.3, 
    -10.46, -10.32, -10.325, -10.44, -10.57, -10.73, -10.81, -10.83, -10.85, 
    -10.68, -10.515, -10.485, -10.46, -10.375, -10.2, -9.87, -9.71, -9.97, 
    -10.115, -10.29, -10.265, -10.525, -10.655, -10.83, -11.13, -11.32, 
    -11.45, -11.365, -11.41, -11.175, -11, -11.05, -11.16, -11.21, -11.25, 
    -11.325, -11.46, -11.74, -11.78, -11.23, -10.245, -9.775, -9.115, -8.925, 
    -10.265, -10.64, -11.025, -11.22, -11.205, -11.165, -11, -10.64, -10.21, 
    -9.67, -8.725, -7.44, -7.26, -7.165, -6.45, -6.07, -5.98, -5.965, -5.635, 
    -4.63, -3.835, -3.85, -3.82, -4.06, -3.585, -4.02, -4.765, -5.095, -5.26, 
    -5.36, -5, -4.545, -4.355, -4.075, -4.35, -4.48, -4.435, -4.39, -4.57, 
    -4.73, -5.175, -5.51, -6.235, -6.595, -6.35, -6.12, -6.375, -5.735, 
    -6.26, -6.19, -6.82, -7.175, -7.385, -7.775, -8.295, -8.16, -8.425, 
    -8.16, -7.82, -7.76, -7.835, -7.975, -8.065, -8.135, -8.09, -7.875, 
    -7.91, -7.56, -6.925, -5.675, -5.265, -4.71, -4.275, -5.165, -7.075, 
    -7.53, -8.385, -10.07, -11.04, -9.97, -9.465, -9.525, -9.72, -9.175, 
    -8.805, -9.18, -8.68, -9.065, -9.46, -9.745, -8.465, -6.73, -3.945, 
    -0.485, -0.495, -0.645, -2.17, -4.61, -5.76, -6.04, -6.25, -6.28, -5.96, 
    -6.185, -5.615, -5.485, -5.62, -5.33, -5.25, -5.07, -4.695, -4.665, 
    -4.62, -4.345, -4.385, -4.2, -4.09, -4.535, -3.27, -3.08, -3.26, -3.99, 
    -4.615, -5.075, -5.045, -4.375, -4.35, -4.355, -4.49, -4.785, -4.645, 
    -4.725, -4.53, -4.265, -4.075, -3.99, -3.95, -3.695, -3.64, -3.775, 
    -3.84, -3.81, -3.76, -3.865, -4.39, -4.74, -5.52, -6.44, -7.42, -7.99, 
    -8.725, -10.68, -12.035, -12.77, -12.49, -13.635, -15.155, -15.77, 
    -16.06, -16.15, -15.66, -15.92, -15.74, -12.88, -9.905, -6.055, -4.78, 
    -5.285, -5.765, -7.07, -8.32, -10.375, -12.445, -12.86, -12.95, -13.015, 
    -12.6, -12.31, -11.595, -11.38, -11.495, -11.11, -11.01, -10.505, -10.46, 
    -10.64, -10.375, -7.355, -3.06, -0.025, 0.585, -1.085, -1.615, -2.14, 
    -2.935, -4.09, -4.345, -5.01, -4.615, -4.715, -4.73, -4.525, -4.585, 
    -4.71, -5.085, -4.83, -4.06, -4.135, -4.375, -4.645, -5.415, -4.645, 
    -2.545, -1.125, -0.895, -0.94, -1.635, -2.395, -2.705, -3.54, -4.98, 
    -4.475, -4.38, -4.09, -5.535, -5.845, -5.85, -4.81, -4.02, -4.13, -4.63, 
    -5.645, -5.195, -5.64, -5.865, -2.765, 0.66, 1.53, 1.22, 1.9, 1.68, 1.07, 
    -0.37, -1.655, -3.4, -4.36, -4.665, -4.765, -4.8, -4.94, -5.55, -5.315, 
    -5.13, -4.915, -5.165, -5.695, -5.65, -5.645, -5.63, -1.34, 2.43, 3.78, 
    4.19, 3.38, 3.8, 3.395, 1.47, 0.345, -0.085, -0.675, -0.12, -2.305, 
    -4.25, -4.78, -4.225, -4.34, -5.215, -5.575, -2.12, -3.445, -1.35, 
    -0.435, -0.095, 1.43, 1.76, 2.09, 2.54, 2.19, 1.905, 1.185, 1.175, 
    -0.655, -1.435, -2.045, -1.88, -3.135, -3.9, -3.785, -2.76, -2.755, 
    -2.575, -3.11, -4.3, -5.945, -6.455, -6.14, -5.77, -3.155, 0.405, 2.715, 
    2.23, 2.61, 0.42, 1.26, -0.115, -1.685, -2.155, -2.805, -3.24, -3.125, 
    -3.45, -4.3, -4.965, -5.03, -5.665, -5.7, -5.585, -5.795, -5.925, -6.055, 
    -6.155, -5.78, -5.09, -5.12, -4.5, -4.32, -4.195, -4.57, -5.32, -6.03, 
    -6.63, -7.41, -8.055, -8.335, -8.65, -8.58, -8.6, -9.29, -10.37, -10.12, 
    -9.49, -8.435, -8.325, -9.545, -7.535, -6.17, -4.84, -3.28, -2.545, 
    -2.07, -1.18, -1.835, -2.55, -2.56, -2.47, -2.72, -2.68, -3.175, -3.03, 
    -2.35, -2.535, -3.365, -3.07, -3.2, -3.105, -4.345, -3.715, -3.79, 
    -3.585, -1.015, 0.52, 2.87, 3.41, 2.845, 1.565, 1.67, 0.03, -2.025, 
    -2.87, -3.785, -3.61, -3.735, -3.275, -2.905, -3.425, -2.73, -3.705, 
    -3.81, -4.375, -5.085, -6.665, -5.465, -4.25, -1.75, 1.065, 0.805, 1.4, 
    2.235, 2.115, 1.685, -0.19, -2.595, -4.095, -4.015, -3.665, -3.205, 
    -3.03, -2.985, -3.485, -4.155, -4.565, -5.53, -5.695, -4.95, -5.59, 
    -5.92, -5.84, -5.445, -4.705, -4.615, -3.24, -3.86, -3.725, -4.13, -4.04, 
    -4.295, -4.435, -4.19, -4.33, -4.815, -5.005, -5.065, -4.825, -4.8, 
    -4.64, -4.24, -4.485, -4.825, -4.995, -5.245, -5.265, -5.22, -5.775, 
    -5.79, -5.325, -4.55, -5.65, -5.77, -5.91, -7.145, -7.855, -9.365, -8.31, 
    -7.795, -7.275, -7.145, -7.52, -7.775, -7.36, -7.85, -8.25, -8.15, -8.14, 
    -8.6, -8.595, -7.36, -5.85, -4.705, -5.065, -5.045, -5.975, -5.795, 
    -5.55, -6.68, -7.605, -8.11, -7.86, -7.685, -7.485, -7.135, -7.315, 
    -7.36, -7.205, -6.965, -6.82, -6.835, -6.99, -6.895, -6.84, -6.525, 
    -6.02, -5.675, -4.24, -4.675, -4.665, -4.695, -5.27, -6.405, -7.235, 
    -7.1, -7.345, -7.725, -7.48, -7.275, -7.79, -7.68, -7.6, -7.385, -6.56, 
    -5.955, -6.11, -6.545, -6.635, -6.515, -6.17, -5.305, -5.655, -6.005, 
    -6.695, -7.035, -7.16, -7.205, -7.37, -7.59, -7.7, -7.82, -8.26, -8.495, 
    -8.565, -8.605, -8.81, -9.19, -9.41, -9.475, -9.51, -9.555, -9.64, -9.5, 
    -9.35, -9.2, -9.22, -9.44, -9.615, -9.78, -9.78, -9.685, -9.65, -9.625, 
    -9.6, -9.625, -9.74, -9.875, -9.965, -10.075, -10.175, -10.23, -10.215, 
    -10.255, -10.31, -10.31, -10.375, -10.22, -9.755, -8.63, -7.215, -8.505, 
    -9.28, -9.46, -10.105, -10.5, -10.91, -11.29, -11.585, -11.655, -11.925, 
    -12.14, -12.165, -11.54, -11.055, -11.17, -11.26, -10.815, -10.49, 
    -10.505, -10.025, -9.39, -9.115, -8.83, -8.345, -6.725, -6.045, -5.165, 
    -5.88, -7.2, -7.63, -7.795, -8.485, -10.6, -11.19, -9.17, -8.75, -9.605, 
    -10.255, -10.735, -10.06, -8.325, -6.455, -6.355, -6.43, -5.34, -3.955, 
    -2.875, -3.755, -3.085, -2.67, -2.3, -3.165, -4.445, -5.105, -5.345, 
    -5.525, -6.06, -6.5, -7.16, -7.35, -7.11, -8.16, -8.68, -8.495, -8.6, 
    -8.165, -7.945, -8.435, -6.715, -4.175, -2.98, -2.245, -2.635, -2.99, 
    -3.59, -4.015, -5.26, -6.64, -6.955, -6.945, -6.925, -6.8, -7.245, -7.65, 
    -8, -8.105, -8.07, -7.99, -8.055, -8.935, -9.44, -9.425, -6.345, -4.485, 
    -3.795, -3.12, -2.88, -2.25, -2.125, -3.3, -5.79, -7.66, -8.255, -8.985, 
    -9.48, -9.625, -10.43, -10.325, -9.5, -10.63, -10.7, -10.325, -10.52, 
    -10.815, -10.675, -10.165, -6.18, -3.14, -1.37, -1.145, -0.9, -0.62, 
    -0.66, -3.105, -4.88, -6.73, -6.945, -7.765, -8.805, -8.975, -8.825, 
    -8.2, -7.88, -9.39, -8.385, -8.9, -7.305, -7.37, -9.75, -9.985, -6.56, 
    -1.025, 1.22, 1.44, 0.785, 0.615, 0.5, -1.65, -3.605, -4.805, -5.71, 
    -5.435, -5.24, -5.53, -5.61, -5.725, -6.06, -6.46, -6.985, -7.275, 
    -7.265, -7.285, -7.25, -7.255, -7.085, -6.685, -6.695, -6.635, -6.77, 
    -6.92, -6.815, -7.225, -7.32, -7.365, -7.32, -7.345, -7.475, -7.72, 
    -7.725, -7.9, -8.01, -8.005, -8.005, -8.155, -8.295, -8.405, -8.615, 
    -8.675, -8.375, -7.33, -6.57, -6.145, -7.515, -6.66, -5.42, -6.335, 
    -7.645, -8.825, -9.915, -11.955, -11.91, -11.31, -10.255, -10.925, 
    -10.965, -10.295, -9.375, -9.245, -9.375, -9.755, -10.95, -10.68, -6.425, 
    -0.755, -0.125, -1.15, -2.785, -3.34, -3.385, -3.89, -4.725, -6.705, 
    -7.995, -7.465, -7.3, -7.64, -9.24, -9.84, -10.31, -9.99, -9.83, -9.6, 
    -9.3, -8.495, -7.625, -6.185, -4.885, -5.4, -4.21, -1.24, -1.065, -1.255, 
    -1.425, -2.215, -3.815, -5.24, -5.98, -5.975, -6.325, -6.35, -6.46, 
    -6.48, -6.93, -7.535, -7.795, -8.035, -8.045, -7.93, -8.735, -8.93, 
    -7.295, -6.155, -6.31, -5.095, -4.445, -5.165, -6.095, -5.32, -6.735, 
    -8.38, -9.31, -9.57, -9.25, -9.895, -9.365, -8.545, -8.21, -7.295, -6.67, 
    -7.195, -6.61, -6.67, -6.725, -6.145, -5.555, -5.355, -4.36, -3.695, 
    -4.14, -4.485, -4.5, -4.57, -4.555, -4.615, -4.52, -4.37, -4.4, -4.33, 
    -4.315, -4.195, -4.16, -4.23, -4.41, -4.47, -4.605, -4.95, -5.225, -4.84, 
    -4, -3.795, -2.98, -1.985, -2.375, -2.63, -2.42, -2.535, -4.08, -6.485, 
    -6.71, -5.935, -6.07, -6.475, -6.465, -6.67, -6.925, -7.095, -7.7, -7.6, 
    -7.435, -7.48, -7.89, -8.11, -8.09, -8, -7.58, -7.225, -6.825, -6.825, 
    -6.71, -6.68, -7.045, -8.085, -8.965, -9.575, -9.685, -9.85, -10.19, 
    -10.47, -11.075, -11.385, -11.22, -12.165, -12.885, -14.19, -14.465, 
    -13.165, -6.15, -5.99, -6.675, -5.78, -4.725, -6.39, -7.43, -8.135, 
    -8.98, -10.35, -10.75, -11.035, -12.695, -13.41, -13.825, -14.255, 
    -14.295, -14.6, -15.105, -13.685, -12.32, -11.06, -11.32, -10.655, -9.62, 
    -9.305, -8.37, -8.195, -6.635, -8.045, -7.84, -7.43, -8.675, -11.25, 
    -13.195, -11.835, -12.225, -12.505, -11.32, -11.215, -10.7, -10.465, 
    -10.26, -9.855, -9.795, -9.725, -9.865, -9.715, -8.72, -8.1, -7.4, -6.72, 
    -6.94, -8.03, -7.95, -7.94, -8.505, -8.735, -8.84, -8.865, -9.165, -9.31, 
    -9.26, -9.06, -9.1, -9.045, -8.615, -8.56, -8.64, -8.805, -8.88, -8.76, 
    -8.4, -7.845, -7.49, -7.125, -7.01, -6.955, -6.95, -6.745, -6.995, -7.18, 
    -7.28, -7.07, -7.095, -7.025, -6.625, -6.395, -6.305, -6.3, -6.215, 
    -6.22, -6.33, -6.355, -6.22, -5.985, -5.475, -5.3, -5.195, -4.985, -4.92, 
    -4.855, -5.115, -5.4, -5.455, -5.76, -5.695, -5.47, -5.305, -5.165, 
    -5.085, -5.23, -5.325, -5.285, -5.295, -5.315, -5.375, -5.275, -5.255, 
    -5.175, -4.885, -4.745, -4.825, -4.745, -4.745, -4.535, -5.295, -5.79, 
    -6.865, -8.16, -8.745, -9.715, -10.79, -9.655, -10.88,
  -7.355, -7.545, -6.75, -6.6, -6.515, -6.545, -7.34, -7.17, -5.715, -3.385, 
    -2.5, -2.31, -2.12, -1.97, -1.89, -2.04, -2.135, -3.33, -4.08, -4.8, 
    -5.035, -5.04, -4.9, -5.815, -5.1, -5.15, -5.315, -5.8, -6.785, -6.35, 
    -5.995, -4.845, -0.33, 1.05, 2.065, 2.82, 3.24, 4.18, 5.065, 4.925, 
    3.445, 2.475, 0.415, -2.325, -2.92, -3.28, -3.53, -2.68, -1.465, -2.74, 
    -1.81, -1.145, -0.18, -0.495, -0.52, 0.235, 1.205, 2.535, 2.73, 3.665, 
    4.295, 4.175, 4.94, 4.9, 4.45, 4.64, 2.975, 2.725, 2.615, 2.685, 2.435, 
    1.81, 0.91, 0.205, -0.235, -0.47, -0.515, -0.64, -0.845, -1.78, -2.05, 
    -1.92, -2.125, -1.23, -1.25, -1.145, -1.6, -1.23, -1.585, -1.585, -2.3, 
    -3.15, -3.33, -3.36, -3.455, -3.855, -4.075, -4.75, -4.96, -5.165, 
    -5.515, -5.835, -6.545, -6.57, -5.72, -5.005, -4.595, -4.815, -3.385, 
    -3.49, -4.83, -4.685, -4.665, -4.815, -4.99, -5.62, -5.855, -6.195, 
    -6.57, -7.72, -6.98, -8.075, -8.33, -7.45, -7.99, -9.205, -9.06, -7.505, 
    -3.675, -0.52, -1.075, 0.005, 0.47, 0.59, 1.325, 1.63, 1.59, -0.02, 
    -1.915, -3.25, -3.25, -2.425, -4.04, -5.65, -5.835, -5.745, -5.095, 
    -5.94, -6.22, -4.83, -5.01, -4.02, 1.03, 3.93, 4.6, 4.285, 5.385, 5.39, 
    5.855, 5.045, 3.88, 2.25, -0.07, -1.25, -1.275, -1.83, -2.23, -2.965, 
    -3.6, -4.115, -3.435, -3.18, -3.76, -4.225, -3.655, -3.03, -2.51, -2.165, 
    0.25, 0.005, 0.1, -0.37, -0.09, 0.575, -0.515, -1.49, -1.795, -1.965, 
    -2.835, -2.945, -2.88, -3.1, -3.305, -3.18, -3.02, -3.015, -2.87, -2.635, 
    -2.615, -2.5, -2.25, -1.475, -1.045, -0.975, -0.885, -0.44, 0.04, 0.575, 
    0.585, 0.22, -0.6, -1.41, -1.905, -2.355, -2.885, -3.295, -3.56, -3.7, 
    -3.8, -4.255, -4.765, -5.17, -5.03, -5.185, -4.64, -3.875, -3.515, 
    -1.445, -0.825, -1.09, -1.695, -2.995, -3.1, -3.2, -3.325, -3.35, -3.39, 
    -3.75, -3.445, -3.285, -3.715, -4.055, -3.645, -3.545, -3.24, -2.81, 
    -2.575, -2.42, -2.11, -1.765, -1.535, -1.51, -1.54, -1.775, -1.7, -0.625, 
    -0.39, -0.87, -1.65, -2.055, -2.42, -2.41, -2.55, -2.84, -2.545, -2.04, 
    -2.205, -2.17, -2.405, -3.215, -3.525, -3.61, 0.655, 3.6, 5.785, 6.57, 
    6.995, 7.15, 7.53, 7.385, 5.8, 4.335, 4.11, 4.4, 4.24, 4.335, 4.73, 
    4.535, 2.89, 1.555, 0.325, 0.35, 0.845, 0.995, 0.935, 1.355, 1.905, 
    4.155, 4.245, 4.125, 6.345, 5.6, 5.915, 5.98, 5.43, 4.75, 4.135, 3.435, 
    1.83, 1.76, 2.32, 1.64, 0.425, 0.01, -0.145, -0.32, -0.23, -0.18, -0.03, 
    0.285, 0.6, 1.02, 1.555, 2.43, 3, 4.035, 3.705, 3.68, 3.845, 3.64, 2.905, 
    3.01, 3.07, 3.265, 3.21, 2.86, 2.855, 2.865, 2.67, 2.83, 2.345, 1.865, 
    1.64, 1.73, 3.605, 3.61, 3.465, 3.61, 4.065, 4.53, 5.265, 5.195, 5.21, 
    4.105, 3.33, 3.12, 2.525, 1.895, 0.15, 1.09, 0, -0.015, -0.63, 0.365, 
    0.835, -0.315, -0.39, -0.23, 4.315, 6.37, 6.895, 7.54, 8.86, 9.645, 
    9.965, 10.18, 9.68, 7.155, 4.065, 3.22, 3.015, 2.745, 2.37, 2.38, 2.035, 
    2.295, 1.67, 3.37, 4.295, 3.935, 3.145, 3.32, 8.21, 11.115, 11.675, 
    12.655, 13.19, 13.435, 13.86, 13.49, 12.665, 10.17, 7.065, 5.96, 5.635, 
    5.365, 5.86, 5.51, 6.28, 7.3, 6.65, 6.65, 6.48, 6.695, 5.76, 5.82, 10.15, 
    11.875, 13.14, 14.395, 14.8, 14.755, 14.34, 14.805, 13.355, 10.935, 
    8.645, 7.925, 8.335, 8.8, 9.5, 9.395, 9.405, 9.295, 9.275, 8.95, 8.11, 
    6.99, 5.58, 2.68, 3.73, 6.09, 8.08, 7.55, 8.205, 8.445, 7.735, 7.105, 
    3.555, 1.365, 1.605, 0.555, -0.095, -0.245, -0.26, -0.435, -0.365, 
    -0.355, -0.08, -0.255, -0.205, -0.09, -0.065, -0.125, -0.135, 0.01, 
    1.385, 1.325, 2.04, 1.44, 0.56, 1.59, 2, 0.745, -0.065, -1.02, -1.85, 
    -2.13, -2.685, -2.695, -2.875, -2.955, -3.25, -3.665, -3.755, -3.6, 
    -3.76, -3.7, -0.905, -0.065, 1.235, 1.45, 1.37, 1.02, 2.045, 3.05, 2.44, 
    0.715, 0.185, -0.005, -0.605, -0.89, -0.365, -0.47, -0.855, -0.65, 
    -0.475, -0.29, -0.12, -0.145, -1.565, -1.24, -0.695, 0.885, 3.405, 3.905, 
    4.145, 5.08, 5.135, 4.29, 3.015, 1.875, 1.085, 0.55, 0.14, -0.35, -0.775, 
    -1.04, -1.3, -1.82, -2.17, -1.585, -2.265, -1.475, -1.1, -0.55, -0.065, 
    0.42, 1.105, 1.775, 1.865, 1.84, 1.32, 1.39, 1.325, 1.255, 0.875, 1.505, 
    1.655, 0.38, -0.1, -0.275, -0.385, -0.22, 0.45, 0.43, 0.49, 0.57, 0.58, 
    0.53, 0.44, 0.31, 0.385, 0.665, 1.135, 0.99, 1.275, 0.67, 0.04, -1.21, 
    -2.36, -3.435, -3.77, -4.13, -4.62, -4.36, -5.16, -5.175, -5.795, -6.895, 
    -7.15, -7.68, -8.83, -8.525, -5.37, -3.675, -2.575, -2.4, -1.495, -1.24, 
    -1.025, -0.9, -1.645, -3.29, -4.665, -5.31, -6.23, -6.83, -6.85, -6.555, 
    -6.935, -6.27, -5.78, -4.76, -4.385, -5.055, -4.825, -4.195, -2.995, 
    -0.53, 0.425, 0.46, 1.77, 2.12, 1.37, 1.625, 0.675, -0.295, -0.265, 0.47, 
    0.575, 0.845, 1.185, 2.2, 1.26, -1.705, -3.45, -4.61, -5.7, -7.2, -7.61, 
    -7.88, -8.115, -8.325, -8.22, -6.61, -5.275, -5.45, -5.67, -7.43, -8.115, 
    -9.05, -9.905, -9.425, -9.425, -9.975, -10.41, -10.37, -10.525, -10.585, 
    -10.59, -10.185, -10.37, -10.9, -10.375, -10.3, -9.47, -7.345, -4.955, 
    -4.905, -4.81, -3.835, -3.385, -4.11, -4.87, -6.115, -6.84, -7.425, 
    -7.925, -8.435, -8.58, -8.355, -8.895, -9.32, -10.21, -11.555, -10.74, 
    -9.74, -11.12, -11.795, -8.96, -8.105, -6.325, -5.97, -5.05, -4.475, 
    -5.55, -6.345, -7.165, -8.095, -8.82, -9.12, -9.48, -9.46, -9.425, 
    -9.385, -9.26, -8.82, -8.485, -8.135, -7.27, -6.12, -5.78, -4.615, 
    -3.995, -4.02, -4.47, -3.84, -3.655, -3.445, -2.9, -2.355, -2.185, 
    -2.095, -1.985, -1.8, -1.595, -1.53, -1.515, -1.49, -1.565, -1.435, 
    -1.435, -1.68, -1.955, -2.365, -2.435, -2.37, -1.365, -0.055, 0.575, 1.5, 
    3.035, 3.68, 4.335, 4.95, 3.63, 1.775, 0.865, 0.36, 0.275, 0.995, 1.82, 
    1.785, 1.4, 1.36, 1.285, 1.6, 1.835, 1.875, 1.515, 1.73, 3.245, 4.875, 
    5.565, 6.04, 5.82, 5.32, 5.02, 4.055, 4.01, 3.235, 2.145, 1.935, 1.62, 
    1.66, 1.345, 1.35, 0.745, 0.8, 0.725, 0.695, 0.09, 0.1, -0.44, -0.665, 
    1.735, 4.885, 5.61, 6.485, 6.69, 6.055, 6.27, 5.845, 5.125, 3.245, 1.01, 
    0.41, 1.095, 0.325, 0.5, 0.305, 0.655, 1.325, 1.02, 1.255, 0.355, 0.56, 
    0.72, 0.96, 3.15, 5.19, 5.59, 7.01, 7.335, 7.925, 7.875, 7.895, 6.835, 
    4.98, 2.54, 0.655, 0.6, 0.4, 0.27, 0.49, 0.76, 0.82, 1.415, 3.575, 4.175, 
    1.61, 1.81, 1.805, 5.895, 10.93, 11.875, 12.64, 13.65, 14.125, 14.33, 
    13.455, 11.69, 8.375, 6.52, 6.475, 8.25, 8.96, 7.66, 7.7, 7.52, 7.625, 
    7.815, 6.98, 4.965, 3.055, 2.155, 4.905, 7.49, 9.84, 11.135, 12.03, 
    12.36, 11.785, 12.515, 10.92, 10.01, 8.255, 7.295, 6.835, 7.165, 7.89, 
    8.21, 7.47, 6.67, 6.075, 6.055, 5.65, 5.05, 4.79, 4.53, 4.405, 4.635, 
    6.24, 6.61, 6.805, 7.015, 6.83, 6.02, 4.875, 4.105, 3.2, 2.305, 2.36, 
    2.155, 1.6, 1.145, 0.875, 0.415, -0.01, -0.35, -0.21, -0.37, -0.445, 
    -0.4, -0.04, 0.475, 2.315, 3.425, 4.885, 5.01, 3.305, 2.65, 1.91, 2.11, 
    1.01, -0.785, -2.23, -2.46, -2.97, -3.2, -2.71, -2.51, -2.93, -3.775, 
    -4.095, -4.535, -4.84, -6.07, -6.715, -3.515, -0.39, -0.05, -0.225, 0.32, 
    0.97, 1.155, 0.89, 0.04, -2.045, -3.91, -4.535, -4.6, -5.05, -5.16, 
    -4.72, -4.505, -5.255, -6.435, -6.42, -5.605, -5.01, -5.03, -4.77, 
    -2.195, 2.48, 4.08, 5.16, 5.565, 5.865, 6.11, 5.7, 4.06, 1.125, 0.435, 
    1.28, 0.965, 0.3, 1.215, 0.53, 0.51, 1.36, 0.055, -0.23, -0.62, 0, 0.895, 
    0.905, 1.045, 2.225, 3.185, 4.6, 4.88, 5.415, 4.655, 4.425, 3.8, 1.905, 
    -0.445, -1.38, -1.93, -1.92, 0.985, 2.22, 2.435, 1.735, 1.81, 2.32, 
    2.415, 1.915, 0.91, 2.285, 2.85, 5.575, 7.23, 8.69, 8.46, 7.6, 6.61, 6.31, 
    6.02, 5.235, 4.925, 4.94, 4.37, 3.765, 5.105, 5.15, 4.895, 4.455, 3.955, 
    3.905, 3.905, 3.665, 3.23, 2.34, 2.375, 2.05, 0.97, 0.635, -1.855, -2.95, 
    -3.085, -3.63, -4.23, -5.015, -5.825, -6.425, -7.33, -8.405, -8.91, 
    -8.615, -9.645, -10.04, -10.88, -11.45, -11.965, -12.235, -12.515, 
    -12.415, -10.93, -8.25, -6.695, -6.955, -5.96, -7.365, -6.795, -7.075, 
    -7.945, -9.305, -11.035, -11.44, -11.825, -11.58, -12.035, -12.755, 
    -12.61, -11.075, -10.5, -10.245, -9.655, -9.535, -9.825, -9.65, -9.095, 
    -8.31, -7.095, -7.035, -6.855, -7.495, -8.515, -9.36, -9.965, -10.825, 
    -11.33, -11.56, -11.925, -12.32, -12.825, -12.88, -13.815, -14.32, 
    -14.955, -14.53, -14.415, -14.87, -14.375, -14.77, -14.145, -10.085, 
    -9.09, -8.33, -6.735, -7.955, -7.56, -8.015, -9.275, -10.56, -12.09, 
    -12.675, -13.005, -12.425, -11.535, -10.825, -10.895, -10.755, -10.785, 
    -10.695, -10.23, -10.43, -10.04, -9.725, -7.485, -1.285, -0.29, -0.16, 
    -0.38, -0.045, -0.255, 0.37, -1.49, -2.965, -3.435, -3.87, -3.155, 
    -2.305, -2.33, -2.59, -2.8, -1.925, -1.735, -1.4, -2.195, -2.29, -0.96, 
    -2.005, 0.03, 5.11, 6.15, 6.175, 7.57, 7.14, 7.885, 6.83, 4.14, 0.645, 
    -0.96, -0.375, -0.04, -0.23, -0.145, -0.28, -1.02, 0.615, 0.77, 0.62, 
    0.16, 0.315, -0.91, -2.27, -0.615, 4.14, 4.54, 3.83, 3.195, 3.43, 3.36, 
    2.745, 0.845, -0.315, -1.91, -2.33, -2.745, -3.535, -4.07, -5.01, -5.47, 
    -5.905, -7.04, -7.385, -7.685, -7.2, -6.375, -6.535, -5.69, -3.28, 
    -0.525, 0.79, 0.905, 1.02, 1.56, 1.49, -0.495, -2.175, -2.895, -3.095, 
    -3.4, -2.645, -1.965, -2.055, -2.165, -2.97, -4.335, -3.815, -2.18, 0.21, 
    0.665, 0.43, 0.655, 3.58, 3.495, 4.245, 4.465, 4.85, 4.59, 4.26, 3.67, 
    2.045, 1.785, 2.055, 2.625, 2.445, 2.395, 2.105, 1.475, 0.92, -0.795, 
    -2.14, -3.39, -5.35, -5.66, -5.84, -6.37, -6.355, -6.04, -6.16, -6.745, 
    -6.245, -6.955, -7.37, -8, -8.72, -9.125, -9.62, -10.505, -11.24, -11.81, 
    -12.43, -12.6, -13.06, -13.38, -11.865, -10.825, -10.53, -11.27, -10.905, 
    -9.55, -7.595, -4.085, -3.155, -4.43, -5.375, -6.38, -6.51, -6.2, -7.65, 
    -8.285, -8.77, -9.165, -9.735, -10.02, -10.195, -10.51, -10.71, -10.93, 
    -11.065, -11, -11.06, -11.17, -11.32, -11.375, -10.61, -9.92, -8.895, 
    -8.965, -8.75, -8.755, -9.17, -10.595, -10.675, -10.62, -11.175, -11.345, 
    -11.39, -11.695, -11.66, -11.335, -11.495, -12.24, -12.115, -12.18, 
    -12.14, -11.995, -11.935, -10.885, -7.475, -4.39, -2.31, -2.73, -2.565, 
    -1.045, -1.31, -3.53, -4.64, -4.62, -4.335, -5.515, -5.86, -5.425, 
    -5.865, -5.865, -5.38, -5.42, -5.465, -5.11, -4.655, -5, -5.305, -3.68, 
    0.3, 1.87, 2.7, 3.505, 3.69, 4.08, 3.49, 1.735, -0.97, -2.08, -2.675, 
    -3.06, -3.27, -3.89, -3.07, -1.875, -2.305, -2.15, -2.1, -2.715, -2.985, 
    -0.955, -0.215, 0.515, 5.195, 8.785, 9.225, 8.35, 8.725, 7.705, 6.05, 
    3.71, 0.975, -1.16, -2.095, -1.58, -1.835, -0.91, -0.03, -1.605, -1.17, 
    -1.895, -1.175, -1.545, -2.025, -3.73, -3.86, -3.345, 2.315, 3.785, 
    5.015, 4.19, 3.585, 3.145, 2.52, 1.955, -1.575, -3.39, -3.575, -3.205, 
    -2.665, -2.745, -2.525, -2.835, -2.58, -2.665, -2.57, -3.01, -3.335, 
    -3.565, -3.855, -3.535, -2.955, -1.765, 0.75, 1.5, 1.08, 0.455, 0.315, 
    -1.165, -2.665, -3.43, -4.005, -4.715, -5.455, -5.78, -6.79, -7.465, 
    -7.335, -7.735, -7.89, -6.925, -6.36, -5.835, -6.605, -6.105, -2.23, 
    -0.71, 0.665, 1.175, 1.4, 1.33, 0.61, -1.795, -3.185, -4.505, -5.175, 
    -5.71, -6.015, -5.5, -5.5, -5.585, -5.24, -4.56, -4.76, -4.69, -4.35, 
    -4.465, -4.26, -3.565, 1.83, 3.505, 2.76, 2.385, 2.26, 2.495, 1.51, 
    0.325, -1.195, -1.64, -2.145, -2.565, -3.025, -3.54, -3.24, -3.705, 
    -4.01, -4.6, -4.815, -4.81, -4.86, -5.15, -5.755, -5.32, -3.705, -2.425, 
    -1.77, -2.05, -3.41, -4.075, -4.72, -5.075, -5.605, -6.04, -6.7, -7.5, 
    -7.795, -8.12, -8.675, -10.235, -11.22, -11.485, -12.015, -12.63, -13.78, 
    -15.085, -15.58, -14.845, -11.125, -8.695, -6.685, -6.2, -6.495, -6.385, 
    -7.42, -9.66, -11.865, -13.28, -14.14, -14.65, -15.61, -16.54, -16.78, 
    -17.69, -17.96, -18.28, -18.675, -19.345, -19.56, -19.125, -19.805, 
    -19.305, -14.49, -11.81, -11.34, -11.38, -10.775, -10.575, -10.95, 
    -12.405, -14.26, -15.32, -16.83, -15.885, -16.525, -16.755, -16.51, 
    -15.7, -15.335, -15.35, -15.14, -14.785, -14.17, -13.585, -13.835, 
    -14.24, -12.725, -10.805, -9.535, -7.9, -7.18, -6.33, -7.795, -9.215, 
    -10.115, -9.975, -9.47, -9.36, -9.225, -8.995, -9.485, -9.485, -9.63, 
    -10.185, -11.245, -9.905, -9.77, -10.84, -12.165, -12.645, -12.71, 
    -12.485, -11.98, -10.905, -10.755, -11.565, -12.84, -14.165, -15.435, 
    -15.755, -15.655, -16.355, -17.17, -16.77, -16.02, -15.865, -16.38, 
    -17.825, -18.595, -19.02, -19.315, -19.555, -19.755, -19.985, -19.705, 
    -19.19, -18.81, -18.725, -18.26, -18.495, -18.97, -19.66, -20.705, 
    -21.335, -21.745, -22.295, -23.25, -24.245, -24.665, -24.505, -24.485, 
    -24.37, -24.205, -23.345, -22.25, -22.24, -22.17, -22.07, -21.72, 
    -18.895, -19.35, -17.555, -14.885, -12.675, -15.025, -18.625, -17.785, 
    -16.245, -17.095, -16.09, -16.875, -17.51, -18.045, -18.28, -18.3, 
    -18.415, -17.535, -16.975, -17.025, -17.1, -17.755, -18.285, -18.105, 
    -18.125, -17.525, -17.12, -17.48, -18.1, -18.54, -19.775, -20.585, 
    -21.17, -21.385, -21.095, -21.08, -21.235, -20.99, -20.805, -20.515, 
    -20.42, -20.185, -20.075, -20.405, -20.71, -21.015, -20.97, -20.575, 
    -20.225, -19.76, -19.475, -19.22, -19.465, -19.27, -19.115, -19.405, 
    -19.44, -19.37, -19.37, -19.395, -19.415, -19.415, -19.275, -19.17, 
    -19.21, -19.08, -18.99, -18.95, -18.815, -19.28, -18.905, -15.135, 
    -12.275, -11.595, -10.325, -10.455, -11.855, -12.435, -14.485, -15.87, 
    -17.055, -16.975, -16.375, -16.115, -16.07, -16, -15.48, -15.11, -14.535, 
    -14.875, -14.745, -14.215, -13.755, -13.425, -12.825, -10.51, -7.39, 
    -5.575, -4.445, -4.69, -4.975, -6.65, -7.895, -9.725, -11.065, -10.655, 
    -11.37, -10.1, -9.975, -9.885, -9.42, -9.41, -8.945, -8.61, -8.47, 
    -8.175, -7.835, -7.43, -7.385, -7.315, -6.92, -6.52, -6.23, -5.77, -5.79, 
    -6.225, -6.285, -6.125, -5.98, -5.755, -5.645, -5.51, -5.42, -5.425, 
    -5.535, -5.615, -5.5, -5.315, -5.195, -5.08, -5.12, -5.225, -5.365, 
    -5.59, -5.365, -5.44, -5.41, -5.505, -5.91, -6.135, -6.27, -6.38, -6.515, 
    -6.58, -6.55, -6.56, -6.645, -6.965, -7.265, -7.38, -7.825, -7.89, -7.78, 
    -7.7, -7.755, -7.95, -8.075, -8.12, -8.325, -8.255, -7.81, -8.43, -8.73, 
    -8.65, -9.255, -9.505, -9.465, -9.515, -9.92, -10.06, -10.07, -10.025, 
    -9.935, -9.81, -9.62, -8.785, -8.325, -8.485, -8.735, -8.785, -8.92, 
    -5.815, -4.445, -2.155, -2.13, -4.205, -4.08, -5.545, -6.225, -6.72, 
    -6.51, -6.09, -5.84, -5.775, -5.79, -5.185, -5.145, -4.935, -4.48, -4.06, 
    -3.765, -3.84, -4.545, -4.635, -3.765, -2.795, -2.095, -2.21, -2.855, 
    -3.545, -3.3, -3.06, -2.925, -3.525, -3.695, -3.95, -3.685, -3.495, 
    -3.18, -2.925, -3.41, -3.555, -3.325, -3.215, -3.42, -3.67, -3.945, 
    -4.09, -4.305, -4.125, -3.16, -3.65, -3.36, -2.73, -2.61, -3.21, -4.645, 
    -5.35, -5.675, -5.55, -5.51, -5.575, -5.635, -6.055, -6.94, -7.69, 
    -8.405, -9.185, -8.205, -7.705, -7.895, -7.725, -7.58, -6.49, -3.005, 
    -4.335, -3.93, -4.2, -3.965, -5.115, -6.095, -7.21, -7.88, -8.145, 
    -8.285, -8.885, -8.875, -8.96, -9.115, -8.93, -9.305, -9.47, -9.33, 
    -7.835, -7.315, -7.565, -7.18, -6.55, -5.3, -4.76, -4.48, -4.66, -4.61, 
    -4.58, -4.835, -5.255, -5.445, -5.325, -5.35, -5.245, -5.005, -4.79, 
    -4.74, -4.655, -4.06, -3.845, -3.125, -3.29, -2.995, -3.185, -3.31, 
    -2.025, 1.175, 2.505, 3.175, 3.145, 2.57, 1.095, -1.35, -2.875, -3.63, 
    -4.415, -5.305, -5.74, -4.94, -4.63, -4.425, -4.875, -5.035, -4.79, 
    -5.865, -5.805, -5.955, -5.34, -5.38, -2.91, -0.385, -0.27, 0.215, -0.42, 
    -0.215, -1.255, -2.87, -4.465, -5.465, -7.125, -7.495, -6.945, -5.57, 
    -5.24, -4.35, -4.25, -4.575, -4.62, -4.525, -4.58, -5.09, -5.075, -5.31, 
    -5.065, -4.22, -4.815, -5.265, -5.525, -6.25, -6.02, -6.115, -6.55, 
    -6.92, -6.215, -5.89, -5.82, -5.755, -5.795, -6.735, -8.43, -9.43, -8.76, 
    -8.13, -7.59, -7.745, -8.195, -8.035, -7.89, -7.93, -8.515, -8.45, -8.89, 
    -9.35, -10.29, -11.62, -12.92, -13.94, -14.675, -15.21, -16, -16.61, 
    -16.38, -17.19, -17.32, -17.855, -17.57, -18.915, -18.505, -17.815, 
    -18.93, -19.07, -15.53, -13.015, -12.67, -12.56, -12.655, -11.455, 
    -12.965, -14.29, -15.45, -15.815, -15.785, -15.355, -14.63, -14.145, 
    -14.09, -14.285, -14.1, -13.745, -13.875, -14.36, -14.435, -13.25, -12.4, 
    -12.58, -11.29, -8.965, -8.625, -8.975, -9.55, -10.125, -11.08, -11.315, 
    -12.695, -13.315, -13.875, -13.795, -14.37, -14.84, -13.87, -13.465, 
    -13.915, -14.755, -15.205, -15.305, -15.57, -15.355, -15.43, -14.65, 
    -9.12, -4.545, -3, -5.655, -6.365, -6.82, -6.97, -8.125, -10.44, -12.505, 
    -12.785, -12.57, -11.98, -11.945, -12.24, -11.8, -11.285, -10.035, 
    -10.09, -9.615, -10.11, -10.335, -9.92, -10.165, -7.91, -5.725, -5.41, 
    -5.31, -5.18, -5.97, -6.53, -7.595, -8.935, -9.815, -10.375, -10.545, 
    -11.495, -11.895, -12.705, -12.995, -12.85, -13.365, -12.865, -13.145, 
    -13.335, -13.625, -11.99, -12.155, -7.805, -2.85, -2.62, -2.51, -2.495, 
    -2.89, -3.86, -5.75, -8.58, -10.49, -9.89, -9.2, -9.57, -9.025, -9.41, 
    -9.21, -10.37, -10.85, -10.56, -9.405, -9.39, -10.125, -10.545, -9.535, 
    -8.555, -7.765, -8.935, -8.975, -8.225, -8.225, -8.305, -9.36, -10.3, 
    -10.46, -10.32, -10.325, -10.44, -10.57, -10.73, -10.81, -10.83, -10.85, 
    -10.68, -10.515, -10.485, -10.46, -10.375, -10.2, -9.87, -9.71, -9.97, 
    -10.115, -10.29, -10.265, -10.525, -10.655, -10.83, -11.13, -11.32, 
    -11.45, -11.365, -11.41, -11.175, -11, -11.05, -11.16, -11.21, -11.25, 
    -11.325, -11.46, -11.74, -11.78, -11.23, -10.245, -9.775, -9.115, -8.925, 
    -10.265, -10.64, -11.025, -11.22, -11.205, -11.165, -11, -10.64, -10.21, 
    -9.67, -8.725, -7.44, -7.26, -7.165, -6.45, -6.07, -5.98, -5.965, -5.635, 
    -4.63, -3.835, -3.85, -3.82, -4.06, -3.585, -4.02, -4.765, -5.095, -5.26, 
    -5.36, -5, -4.545, -4.355, -4.075, -4.35, -4.48, -4.435, -4.39, -4.57, 
    -4.73, -5.175, -5.51, -6.235, -6.595, -6.35, -6.12, -6.375, -5.735, 
    -6.26, -6.19, -6.82, -7.175, -7.385, -7.775, -8.295, -8.16, -8.425, 
    -8.16, -7.82, -7.76, -7.835, -7.975, -8.065, -8.135, -8.09, -7.875, 
    -7.91, -7.56, -6.925, -5.675, -5.265, -4.71, -4.275, -5.165, -7.075, 
    -7.53, -8.385, -10.07, -11.04, -9.97, -9.465, -9.525, -9.72, -9.175, 
    -8.805, -9.18, -8.68, -9.065, -9.46, -9.745, -8.465, -6.73, -3.945, 
    -0.485, -0.495, -0.645, -2.17, -4.61, -5.76, -6.04, -6.25, -6.28, -5.96, 
    -6.185, -5.615, -5.485, -5.62, -5.33, -5.25, -5.07, -4.695, -4.665, 
    -4.62, -4.345, -4.385, -4.2, -4.09, -4.535, -3.27, -3.08, -3.26, -3.99, 
    -4.615, -5.075, -5.045, -4.375, -4.35, -4.355, -4.49, -4.785, -4.645, 
    -4.725, -4.53, -4.265, -4.075, -3.99, -3.95, -3.695, -3.64, -3.775, 
    -3.84, -3.81, -3.76, -3.865, -4.39, -4.74, -5.52, -6.44, -7.42, -7.99, 
    -8.725, -10.68, -12.035, -12.77, -12.49, -13.635, -15.155, -15.77, 
    -16.06, -16.15, -15.66, -15.92, -15.74, -12.88, -9.905, -6.055, -4.78, 
    -5.285, -5.765, -7.07, -8.32, -10.375, -12.445, -12.86, -12.95, -13.015, 
    -12.6, -12.31, -11.595, -11.38, -11.495, -11.11, -11.01, -10.505, -10.46, 
    -10.64, -10.375, -7.355, -3.06, -0.025, 0.585, -1.085, -1.615, -2.14, 
    -2.935, -4.09, -4.345, -5.01, -4.615, -4.715, -4.73, -4.525, -4.585, 
    -4.71, -5.085, -4.83, -4.06, -4.135, -4.375, -4.645, -5.415, -4.645, 
    -2.545, -1.125, -0.895, -0.94, -1.635, -2.395, -2.705, -3.54, -4.98, 
    -4.475, -4.38, -4.09, -5.535, -5.845, -5.85, -4.81, -4.02, -4.13, -4.63, 
    -5.645, -5.195, -5.64, -5.865, -2.765, 0.66, 1.53, 1.22, 1.9, 1.68, 1.07, 
    -0.37, -1.655, -3.4, -4.36, -4.665, -4.765, -4.8, -4.94, -5.55, -5.315, 
    -5.13, -4.915, -5.165, -5.695, -5.65, -5.645, -5.63, -1.34, 2.43, 3.78, 
    4.19, 3.38, 3.8, 3.395, 1.47, 0.345, -0.085, -0.675, -0.12, -2.305, 
    -4.25, -4.78, -4.225, -4.34, -5.215, -5.575, -2.12, -3.445, -1.35, 
    -0.435, -0.095, 1.43, 1.76, 2.09, 2.54, 2.19, 1.905, 1.185, 1.175, 
    -0.655, -1.435, -2.045, -1.88, -3.135, -3.9, -3.785, -2.76, -2.755, 
    -2.575, -3.11, -4.3, -5.945, -6.455, -6.14, -5.77, -3.155, 0.405, 2.715, 
    2.23, 2.61, 0.42, 1.26, -0.115, -1.685, -2.155, -2.805, -3.24, -3.125, 
    -3.45, -4.3, -4.965, -5.03, -5.665, -5.7, -5.585, -5.795, -5.925, -6.055, 
    -6.155, -5.78, -5.09, -5.12, -4.5, -4.32, -4.195, -4.57, -5.32, -6.03, 
    -6.63, -7.41, -8.055, -8.335, -8.65, -8.58, -8.6, -9.29, -10.37, -10.12, 
    -9.49, -8.435, -8.325, -9.545, -7.535, -6.17, -4.84, -3.28, -2.545, 
    -2.07, -1.18, -1.835, -2.55, -2.56, -2.47, -2.72, -2.68, -3.175, -3.03, 
    -2.35, -2.535, -3.365, -3.07, -3.2, -3.105, -4.345, -3.715, -3.79, 
    -3.585, -1.015, 0.52, 2.87, 3.41, 2.845, 1.565, 1.67, 0.03, -2.025, 
    -2.87, -3.785, -3.61, -3.735, -3.275, -2.905, -3.425, -2.73, -3.705, 
    -3.81, -4.375, -5.085, -6.665, -5.465, -4.25, -1.75, 1.065, 0.805, 1.4, 
    2.235, 2.115, 1.685, -0.19, -2.595, -4.095, -4.015, -3.665, -3.205, 
    -3.03, -2.985, -3.485, -4.155, -4.565, -5.53, -5.695, -4.95, -5.59, 
    -5.92, -5.84, -5.445, -4.705, -4.615, -3.24, -3.86, -3.725, -4.13, -4.04, 
    -4.295, -4.435, -4.19, -4.33, -4.815, -5.005, -5.065, -4.825, -4.8, 
    -4.64, -4.24, -4.485, -4.825, -4.995, -5.245, -5.265, -5.22, -5.775, 
    -5.79, -5.325, -4.55, -5.65, -5.77, -5.91, -7.145, -7.855, -9.365, -8.31, 
    -7.795, -7.275, -7.145, -7.52, -7.775, -7.36, -7.85, -8.25, -8.15, -8.14, 
    -8.6, -8.595, -7.36, -5.85, -4.705, -5.065, -5.045, -5.975, -5.795, 
    -5.55, -6.68, -7.605, -8.11, -7.86, -7.685, -7.485, -7.135, -7.315, 
    -7.36, -7.205, -6.965, -6.82, -6.835, -6.99, -6.895, -6.84, -6.525, 
    -6.02, -5.675, -4.24, -4.675, -4.665, -4.695, -5.27, -6.405, -7.235, 
    -7.1, -7.345, -7.725, -7.48, -7.275, -7.79, -7.68, -7.6, -7.385, -6.56, 
    -5.955, -6.11, -6.545, -6.635, -6.515, -6.17, -5.305, -5.655, -6.005, 
    -6.695, -7.035, -7.16, -7.205, -7.37, -7.59, -7.7, -7.82, -8.26, -8.495, 
    -8.565, -8.605, -8.81, -9.19, -9.41, -9.475, -9.51, -9.555, -9.64, -9.5, 
    -9.35, -9.2, -9.22, -9.44, -9.615, -9.78, -9.78, -9.685, -9.65, -9.625, 
    -9.6, -9.625, -9.74, -9.875, -9.965, -10.075, -10.175, -10.23, -10.215, 
    -10.255, -10.31, -10.31, -10.375, -10.22, -9.755, -8.63, -7.215, -8.505, 
    -9.28, -9.46, -10.105, -10.5, -10.91, -11.29, -11.585, -11.655, -11.925, 
    -12.14, -12.165, -11.54, -11.055, -11.17, -11.26, -10.815, -10.49, 
    -10.505, -10.025, -9.39, -9.115, -8.83, -8.345, -6.725, -6.045, -5.165, 
    -5.88, -7.2, -7.63, -7.795, -8.485, -10.6, -11.19, -9.17, -8.75, -9.605, 
    -10.255, -10.735, -10.06, -8.325, -6.455, -6.355, -6.43, -5.34, -3.955, 
    -2.875, -3.755, -3.085, -2.67, -2.3, -3.165, -4.445, -5.105, -5.345, 
    -5.525, -6.06, -6.5, -7.16, -7.35, -7.11, -8.16, -8.68, -8.495, -8.6, 
    -8.165, -7.945, -8.435, -6.715, -4.175, -2.98, -2.245, -2.635, -2.99, 
    -3.59, -4.015, -5.26, -6.64, -6.955, -6.945, -6.925, -6.8, -7.245, -7.65, 
    -8, -8.105, -8.07, -7.99, -8.055, -8.935, -9.44, -9.425, -6.345, -4.485, 
    -3.795, -3.12, -2.88, -2.25, -2.125, -3.3, -5.79, -7.66, -8.255, -8.985, 
    -9.48, -9.625, -10.43, -10.325, -9.5, -10.63, -10.7, -10.325, -10.52, 
    -10.815, -10.675, -10.165, -6.18, -3.14, -1.37, -1.145, -0.9, -0.62, 
    -0.66, -3.105, -4.88, -6.73, -6.945, -7.765, -8.805, -8.975, -8.825, 
    -8.2, -7.88, -9.39, -8.385, -8.9, -7.305, -7.37, -9.75, -9.985, -6.56, 
    -1.025, 1.22, 1.44, 0.785, 0.615, 0.5, -1.65, -3.605, -4.805, -5.71, 
    -5.435, -5.24, -5.53, -5.61, -5.725, -6.06, -6.46, -6.985, -7.275, 
    -7.265, -7.285, -7.25, -7.255, -7.085, -6.685, -6.695, -6.635, -6.77, 
    -6.92, -6.815, -7.225, -7.32, -7.365, -7.32, -7.345, -7.475, -7.72, 
    -7.725, -7.9, -8.01, -8.005, -8.005, -8.155, -8.295, -8.405, -8.615, 
    -8.675, -8.375, -7.33, -6.57, -6.145, -7.515, -6.66, -5.42, -6.335, 
    -7.645, -8.825, -9.915, -11.955, -11.91, -11.31, -10.255, -10.925, 
    -10.965, -10.295, -9.375, -9.245, -9.375, -9.755, -10.95, -10.68, -6.425, 
    -0.755, -0.125, -1.15, -2.785, -3.34, -3.385, -3.89, -4.725, -6.705, 
    -7.995, -7.465, -7.3, -7.64, -9.24, -9.84, -10.31, -9.99, -9.83, -9.6, 
    -9.3, -8.495, -7.625, -6.185, -4.885, -5.4, -4.21, -1.24, -1.065, -1.255, 
    -1.425, -2.215, -3.815, -5.24, -5.98, -5.975, -6.325, -6.35, -6.46, 
    -6.48, -6.93, -7.535, -7.795, -8.035, -8.045, -7.93, -8.735, -8.93, 
    -7.295, -6.155, -6.31, -5.095, -4.445, -5.165, -6.095, -5.32, -6.735, 
    -8.38, -9.31, -9.57, -9.25, -9.895, -9.365, -8.545, -8.21, -7.295, -6.67, 
    -7.195, -6.61, -6.67, -6.725, -6.145, -5.555, -5.355, -4.36, -3.695, 
    -4.14, -4.485, -4.5, -4.57, -4.555, -4.615, -4.52, -4.37, -4.4, -4.33, 
    -4.315, -4.195, -4.16, -4.23, -4.41, -4.47, -4.605, -4.95, -5.225, -4.84, 
    -4, -3.795, -2.98, -1.985, -2.375, -2.63, -2.42, -2.535, -4.08, -6.485, 
    -6.71, -5.935, -6.07, -6.475, -6.465, -6.67, -6.925, -7.095, -7.7, -7.6, 
    -7.435, -7.48, -7.89, -8.11, -8.09, -8, -7.58, -7.225, -6.825, -6.825, 
    -6.71, -6.68, -7.045, -8.085, -8.965, -9.575, -9.685, -9.85, -10.19, 
    -10.47, -11.075, -11.385, -11.22, -12.165, -12.885, -14.19, -14.465, 
    -13.165, -6.15, -5.99, -6.675, -5.78, -4.725, -6.39, -7.43, -8.135, 
    -8.98, -10.35, -10.75, -11.035, -12.695, -13.41, -13.825, -14.255, 
    -14.295, -14.6, -15.105, -13.685, -12.32, -11.06, -11.32, -10.655, -9.62, 
    -9.305, -8.37, -8.195, -6.635, -8.045, -7.84, -7.43, -8.675, -11.25, 
    -13.195, -11.835, -12.225, -12.505, -11.32, -11.215, -10.7, -10.465, 
    -10.26, -9.855, -9.795, -9.725, -9.865, -9.715, -8.72, -8.1, -7.4, -6.72, 
    -6.94, -8.03, -7.95, -7.94, -8.505, -8.735, -8.84, -8.865, -9.165, -9.31, 
    -9.26, -9.06, -9.1, -9.045, -8.615, -8.56, -8.64, -8.805, -8.88, -8.76, 
    -8.4, -7.845, -7.49, -7.125, -7.01, -6.955, -6.95, -6.745, -6.995, -7.18, 
    -7.28, -7.07, -7.095, -7.025, -6.625, -6.395, -6.305, -6.3, -6.215, 
    -6.22, -6.33, -6.355, -6.22, -5.985, -5.475, -5.3, -5.195, -4.985, -4.92, 
    -4.855, -5.115, -5.4, -5.455, -5.76, -5.695, -5.47, -5.305, -5.165, 
    -5.085, -5.23, -5.325, -5.285, -5.295, -5.315, -5.375, -5.275, -5.255, 
    -5.175, -4.885, -4.745, -4.825, -4.745, -4.745, -4.535, -5.295, -5.79, 
    -6.865, -8.16, -8.745, -9.715, -10.79, -9.655, -10.88,
  -7.355, -7.545, -6.75, -6.6, -6.515, -6.545, -7.34, -7.17, -5.715, -3.385, 
    -2.5, -2.31, -2.12, -1.97, -1.89, -2.04, -2.135, -3.33, -4.08, -4.8, 
    -5.035, -5.04, -4.9, -5.815, -5.1, -5.15, -5.315, -5.8, -6.785, -6.35, 
    -5.995, -4.845, -0.33, 1.05, 2.065, 2.82, 3.24, 4.18, 5.065, 4.925, 
    3.445, 2.475, 0.415, -2.325, -2.92, -3.28, -3.53, -2.68, -1.465, -2.74, 
    -1.81, -1.145, -0.18, -0.495, -0.52, 0.235, 1.205, 2.535, 2.73, 3.665, 
    4.295, 4.175, 4.94, 4.9, 4.45, 4.64, 2.975, 2.725, 2.615, 2.685, 2.435, 
    1.81, 0.91, 0.205, -0.235, -0.47, -0.515, -0.64, -0.845, -1.78, -2.05, 
    -1.92, -2.125, -1.23, -1.25, -1.145, -1.6, -1.23, -1.585, -1.585, -2.3, 
    -3.15, -3.33, -3.36, -3.455, -3.855, -4.075, -4.75, -4.96, -5.165, 
    -5.515, -5.835, -6.545, -6.57, -5.72, -5.005, -4.595, -4.815, -3.385, 
    -3.49, -4.83, -4.685, -4.665, -4.815, -4.99, -5.62, -5.855, -6.195, 
    -6.57, -7.72, -6.98, -8.075, -8.33, -7.45, -7.99, -9.205, -9.06, -7.505, 
    -3.675, -0.52, -1.075, 0.005, 0.47, 0.59, 1.325, 1.63, 1.59, -0.02, 
    -1.915, -3.25, -3.25, -2.425, -4.04, -5.65, -5.835, -5.745, -5.095, 
    -5.94, -6.22, -4.83, -5.01, -4.02, 1.03, 3.93, 4.6, 4.285, 5.385, 5.39, 
    5.855, 5.045, 3.88, 2.25, -0.07, -1.25, -1.275, -1.83, -2.23, -2.965, 
    -3.6, -4.115, -3.435, -3.18, -3.76, -4.225, -3.655, -3.03, -2.51, -2.165, 
    0.25, 0.005, 0.1, -0.37, -0.09, 0.575, -0.515, -1.49, -1.795, -1.965, 
    -2.835, -2.945, -2.88, -3.1, -3.305, -3.18, -3.02, -3.015, -2.87, -2.635, 
    -2.615, -2.5, -2.25, -1.475, -1.045, -0.975, -0.885, -0.44, 0.04, 0.575, 
    0.585, 0.22, -0.6, -1.41, -1.905, -2.355, -2.885, -3.295, -3.56, -3.7, 
    -3.8, -4.255, -4.765, -5.17, -5.03, -5.185, -4.64, -3.875, -3.515, 
    -1.445, -0.825, -1.09, -1.695, -2.995, -3.1, -3.2, -3.325, -3.35, -3.39, 
    -3.75, -3.445, -3.285, -3.715, -4.055, -3.645, -3.545, -3.24, -2.81, 
    -2.575, -2.42, -2.11, -1.765, -1.535, -1.51, -1.54, -1.775, -1.7, -0.625, 
    -0.39, -0.87, -1.65, -2.055, -2.42, -2.41, -2.55, -2.84, -2.545, -2.04, 
    -2.205, -2.17, -2.405, -3.215, -3.525, -3.61, 0.655, 3.6, 5.785, 6.57, 
    6.995, 7.15, 7.53, 7.385, 5.8, 4.335, 4.11, 4.4, 4.24, 4.335, 4.73, 
    4.535, 2.89, 1.555, 0.325, 0.35, 0.845, 0.995, 0.935, 1.355, 1.905, 
    4.155, 4.245, 4.125, 6.345, 5.6, 5.915, 5.98, 5.43, 4.75, 4.135, 3.435, 
    1.83, 1.76, 2.32, 1.64, 0.425, 0.01, -0.145, -0.32, -0.23, -0.18, -0.03, 
    0.285, 0.6, 1.02, 1.555, 2.43, 3, 4.035, 3.705, 3.68, 3.845, 3.64, 2.905, 
    3.01, 3.07, 3.265, 3.21, 2.86, 2.855, 2.865, 2.67, 2.83, 2.345, 1.865, 
    1.64, 1.73, 3.605, 3.61, 3.465, 3.61, 4.065, 4.53, 5.265, 5.195, 5.21, 
    4.105, 3.33, 3.12, 2.525, 1.895, 0.15, 1.09, 0, -0.015, -0.63, 0.365, 
    0.835, -0.315, -0.39, -0.23, 4.315, 6.37, 6.895, 7.54, 8.86, 9.645, 
    9.965, 10.18, 9.68, 7.155, 4.065, 3.22, 3.015, 2.745, 2.37, 2.38, 2.035, 
    2.295, 1.67, 3.37, 4.295, 3.935, 3.145, 3.32, 8.21, 11.115, 11.675, 
    12.655, 13.19, 13.435, 13.86, 13.49, 12.665, 10.17, 7.065, 5.96, 5.635, 
    5.365, 5.86, 5.51, 6.28, 7.3, 6.65, 6.65, 6.48, 6.695, 5.76, 5.82, 10.15, 
    11.875, 13.14, 14.395, 14.8, 14.755, 14.34, 14.805, 13.355, 10.935, 
    8.645, 7.925, 8.335, 8.8, 9.5, 9.395, 9.405, 9.295, 9.275, 8.95, 8.11, 
    6.99, 5.58, 2.68, 3.73, 6.09, 8.08, 7.55, 8.205, 8.445, 7.735, 7.105, 
    3.555, 1.365, 1.605, 0.555, -0.095, -0.245, -0.26, -0.435, -0.365, 
    -0.355, -0.08, -0.255, -0.205, -0.09, -0.065, -0.125, -0.135, 0.01, 
    1.385, 1.325, 2.04, 1.44, 0.56, 1.59, 2, 0.745, -0.065, -1.02, -1.85, 
    -2.13, -2.685, -2.695, -2.875, -2.955, -3.25, -3.665, -3.755, -3.6, 
    -3.76, -3.7, -0.905, -0.065, 1.235, 1.45, 1.37, 1.02, 2.045, 3.05, 2.44, 
    0.715, 0.185, -0.005, -0.605, -0.89, -0.365, -0.47, -0.855, -0.65, 
    -0.475, -0.29, -0.12, -0.145, -1.565, -1.24, -0.695, 0.885, 3.405, 3.905, 
    4.145, 5.08, 5.135, 4.29, 3.015, 1.875, 1.085, 0.55, 0.14, -0.35, -0.775, 
    -1.04, -1.3, -1.82, -2.17, -1.585, -2.265, -1.475, -1.1, -0.55, -0.065, 
    0.42, 1.105, 1.775, 1.865, 1.84, 1.32, 1.39, 1.325, 1.255, 0.875, 1.505, 
    1.655, 0.38, -0.1, -0.275, -0.385, -0.22, 0.45, 0.43, 0.49, 0.57, 0.58, 
    0.53, 0.44, 0.31, 0.385, 0.665, 1.135, 0.99, 1.275, 0.67, 0.04, -1.21, 
    -2.36, -3.435, -3.77, -4.13, -4.62, -4.36, -5.16, -5.175, -5.795, -6.895, 
    -7.15, -7.68, -8.83, -8.525, -5.37, -3.675, -2.575, -2.4, -1.495, -1.24, 
    -1.025, -0.9, -1.645, -3.29, -4.665, -5.31, -6.23, -6.83, -6.85, -6.555, 
    -6.935, -6.27, -5.78, -4.76, -4.385, -5.055, -4.825, -4.195, -2.995, 
    -0.53, 0.425, 0.46, 1.77, 2.12, 1.37, 1.625, 0.675, -0.295, -0.265, 0.47, 
    0.575, 0.845, 1.185, 2.2, 1.26, -1.705, -3.45, -4.61, -5.7, -7.2, -7.61, 
    -7.88, -8.115, -8.325, -8.22, -6.61, -5.275, -5.45, -5.67, -7.43, -8.115, 
    -9.05, -9.905, -9.425, -9.425, -9.975, -10.41, -10.37, -10.525, -10.585, 
    -10.59, -10.185, -10.37, -10.9, -10.375, -10.3, -9.47, -7.345, -4.955, 
    -4.905, -4.81, -3.835, -3.385, -4.11, -4.87, -6.115, -6.84, -7.425, 
    -7.925, -8.435, -8.58, -8.355, -8.895, -9.32, -10.21, -11.555, -10.74, 
    -9.74, -11.12, -11.795, -8.96, -8.105, -6.325, -5.97, -5.05, -4.475, 
    -5.55, -6.345, -7.165, -8.095, -8.82, -9.12, -9.48, -9.46, -9.425, 
    -9.385, -9.26, -8.82, -8.485, -8.135, -7.27, -6.12, -5.78, -4.615, 
    -3.995, -4.02, -4.47, -3.84, -3.655, -3.445, -2.9, -2.355, -2.185, 
    -2.095, -1.985, -1.8, -1.595, -1.53, -1.515, -1.49, -1.565, -1.435, 
    -1.435, -1.68, -1.955, -2.365, -2.435, -2.37, -1.365, -0.055, 0.575, 1.5, 
    3.035, 3.68, 4.335, 4.95, 3.63, 1.775, 0.865, 0.36, 0.275, 0.995, 1.82, 
    1.785, 1.4, 1.36, 1.285, 1.6, 1.835, 1.875, 1.515, 1.73, 3.245, 4.875, 
    5.565, 6.04, 5.82, 5.32, 5.02, 4.055, 4.01, 3.235, 2.145, 1.935, 1.62, 
    1.66, 1.345, 1.35, 0.745, 0.8, 0.725, 0.695, 0.09, 0.1, -0.44, -0.665, 
    1.735, 4.885, 5.61, 6.485, 6.69, 6.055, 6.27, 5.845, 5.125, 3.245, 1.01, 
    0.41, 1.095, 0.325, 0.5, 0.305, 0.655, 1.325, 1.02, 1.255, 0.355, 0.56, 
    0.72, 0.96, 3.15, 5.19, 5.59, 7.01, 7.335, 7.925, 7.875, 7.895, 6.835, 
    4.98, 2.54, 0.655, 0.6, 0.4, 0.27, 0.49, 0.76, 0.82, 1.415, 3.575, 4.175, 
    1.61, 1.81, 1.805, 5.895, 10.93, 11.875, 12.64, 13.65, 14.125, 14.33, 
    13.455, 11.69, 8.375, 6.52, 6.475, 8.25, 8.96, 7.66, 7.7, 7.52, 7.625, 
    7.815, 6.98, 4.965, 3.055, 2.155, 4.905, 7.49, 9.84, 11.135, 12.03, 
    12.36, 11.785, 12.515, 10.92, 10.01, 8.255, 7.295, 6.835, 7.165, 7.89, 
    8.21, 7.47, 6.67, 6.075, 6.055, 5.65, 5.05, 4.79, 4.53, 4.405, 4.635, 
    6.24, 6.61, 6.805, 7.015, 6.83, 6.02, 4.875, 4.105, 3.2, 2.305, 2.36, 
    2.155, 1.6, 1.145, 0.875, 0.415, -0.01, -0.35, -0.21, -0.37, -0.445, 
    -0.4, -0.04, 0.475, 2.315, 3.425, 4.885, 5.01, 3.305, 2.65, 1.91, 2.11, 
    1.01, -0.785, -2.23, -2.46, -2.97, -3.2, -2.71, -2.51, -2.93, -3.775, 
    -4.095, -4.535, -4.84, -6.07, -6.715, -3.515, -0.39, -0.05, -0.225, 0.32, 
    0.97, 1.155, 0.89, 0.04, -2.045, -3.91, -4.535, -4.6, -5.05, -5.16, 
    -4.72, -4.505, -5.255, -6.435, -6.42, -5.605, -5.01, -5.03, -4.77, 
    -2.195, 2.48, 4.08, 5.16, 5.565, 5.865, 6.11, 5.7, 4.06, 1.125, 0.435, 
    1.28, 0.965, 0.3, 1.215, 0.53, 0.51, 1.36, 0.055, -0.23, -0.62, 0, 0.895, 
    0.905, 1.045, 2.225, 3.185, 4.6, 4.88, 5.415, 4.655, 4.425, 3.8, 1.905, 
    -0.445, -1.38, -1.93, -1.92, 0.985, 2.22, 2.435, 1.735, 1.81, 2.32, 
    2.415, 1.915, 0.91, 2.285, 2.85, 5.575, 7.23, 8.69, 8.46, 7.6, 6.61, 6.31, 
    6.02, 5.235, 4.925, 4.94, 4.37, 3.765, 5.105, 5.15, 4.895, 4.455, 3.955, 
    3.905, 3.905, 3.665, 3.23, 2.34, 2.375, 2.05, 0.97, 0.635, -1.855, -2.95, 
    -3.085, -3.63, -4.23, -5.015, -5.825, -6.425, -7.33, -8.405, -8.91, 
    -8.615, -9.645, -10.04, -10.88, -11.45, -11.965, -12.235, -12.515, 
    -12.415, -10.93, -8.25, -6.695, -6.955, -5.96, -7.365, -6.795, -7.075, 
    -7.945, -9.305, -11.035, -11.44, -11.825, -11.58, -12.035, -12.755, 
    -12.61, -11.075, -10.5, -10.245, -9.655, -9.535, -9.825, -9.65, -9.095, 
    -8.31, -7.095, -7.035, -6.855, -7.495, -8.515, -9.36, -9.965, -10.825, 
    -11.33, -11.56, -11.925, -12.32, -12.825, -12.88, -13.815, -14.32, 
    -14.955, -14.53, -14.415, -14.87, -14.375, -14.77, -14.145, -10.085, 
    -9.09, -8.33, -6.735, -7.955, -7.56, -8.015, -9.275, -10.56, -12.09, 
    -12.675, -13.005, -12.425, -11.535, -10.825, -10.895, -10.755, -10.785, 
    -10.695, -10.23, -10.43, -10.04, -9.725, -7.485, -1.285, -0.29, -0.16, 
    -0.38, -0.045, -0.255, 0.37, -1.49, -2.965, -3.435, -3.87, -3.155, 
    -2.305, -2.33, -2.59, -2.8, -1.925, -1.735, -1.4, -2.195, -2.29, -0.96, 
    -2.005, 0.03, 5.11, 6.15, 6.175, 7.57, 7.14, 7.885, 6.83, 4.14, 0.645, 
    -0.96, -0.375, -0.04, -0.23, -0.145, -0.28, -1.02, 0.615, 0.77, 0.62, 
    0.16, 0.315, -0.91, -2.27, -0.615, 4.14, 4.54, 3.83, 3.195, 3.43, 3.36, 
    2.745, 0.845, -0.315, -1.91, -2.33, -2.745, -3.535, -4.07, -5.01, -5.47, 
    -5.905, -7.04, -7.385, -7.685, -7.2, -6.375, -6.535, -5.69, -3.28, 
    -0.525, 0.79, 0.905, 1.02, 1.56, 1.49, -0.495, -2.175, -2.895, -3.095, 
    -3.4, -2.645, -1.965, -2.055, -2.165, -2.97, -4.335, -3.815, -2.18, 0.21, 
    0.665, 0.43, 0.655, 3.58, 3.495, 4.245, 4.465, 4.85, 4.59, 4.26, 3.67, 
    2.045, 1.785, 2.055, 2.625, 2.445, 2.395, 2.105, 1.475, 0.92, -0.795, 
    -2.14, -3.39, -5.35, -5.66, -5.84, -6.37, -6.355, -6.04, -6.16, -6.745, 
    -6.245, -6.955, -7.37, -8, -8.72, -9.125, -9.62, -10.505, -11.24, -11.81, 
    -12.43, -12.6, -13.06, -13.38, -11.865, -10.825, -10.53, -11.27, -10.905, 
    -9.55, -7.595, -4.085, -3.155, -4.43, -5.375, -6.38, -6.51, -6.2, -7.65, 
    -8.285, -8.77, -9.165, -9.735, -10.02, -10.195, -10.51, -10.71, -10.93, 
    -11.065, -11, -11.06, -11.17, -11.32, -11.375, -10.61, -9.92, -8.895, 
    -8.965, -8.75, -8.755, -9.17, -10.595, -10.675, -10.62, -11.175, -11.345, 
    -11.39, -11.695, -11.66, -11.335, -11.495, -12.24, -12.115, -12.18, 
    -12.14, -11.995, -11.935, -10.885, -7.475, -4.39, -2.31, -2.73, -2.565, 
    -1.045, -1.31, -3.53, -4.64, -4.62, -4.335, -5.515, -5.86, -5.425, 
    -5.865, -5.865, -5.38, -5.42, -5.465, -5.11, -4.655, -5, -5.305, -3.68, 
    0.3, 1.87, 2.7, 3.505, 3.69, 4.08, 3.49, 1.735, -0.97, -2.08, -2.675, 
    -3.06, -3.27, -3.89, -3.07, -1.875, -2.305, -2.15, -2.1, -2.715, -2.985, 
    -0.955, -0.215, 0.515, 5.195, 8.785, 9.225, 8.35, 8.725, 7.705, 6.05, 
    3.71, 0.975, -1.16, -2.095, -1.58, -1.835, -0.91, -0.03, -1.605, -1.17, 
    -1.895, -1.175, -1.545, -2.025, -3.73, -3.86, -3.345, 2.315, 3.785, 
    5.015, 4.19, 3.585, 3.145, 2.52, 1.955, -1.575, -3.39, -3.575, -3.205, 
    -2.665, -2.745, -2.525, -2.835, -2.58, -2.665, -2.57, -3.01, -3.335, 
    -3.565, -3.855, -3.535, -2.955, -1.765, 0.75, 1.5, 1.08, 0.455, 0.315, 
    -1.165, -2.665, -3.43, -4.005, -4.715, -5.455, -5.78, -6.79, -7.465, 
    -7.335, -7.735, -7.89, -6.925, -6.36, -5.835, -6.605, -6.105, -2.23, 
    -0.71, 0.665, 1.175, 1.4, 1.33, 0.61, -1.795, -3.185, -4.505, -5.175, 
    -5.71, -6.015, -5.5, -5.5, -5.585, -5.24, -4.56, -4.76, -4.69, -4.35, 
    -4.465, -4.26, -3.565, 1.83, 3.505, 2.76, 2.385, 2.26, 2.495, 1.51, 
    0.325, -1.195, -1.64, -2.145, -2.565, -3.025, -3.54, -3.24, -3.705, 
    -4.01, -4.6, -4.815, -4.81, -4.86, -5.15, -5.755, -5.32, -3.705, -2.425, 
    -1.77, -2.05, -3.41, -4.075, -4.72, -5.075, -5.605, -6.04, -6.7, -7.5, 
    -7.795, -8.12, -8.675, -10.235, -11.22, -11.485, -12.015, -12.63, -13.78, 
    -15.085, -15.58, -14.845, -11.125, -8.695, -6.685, -6.2, -6.495, -6.385, 
    -7.42, -9.66, -11.865, -13.28, -14.14, -14.65, -15.61, -16.54, -16.78, 
    -17.69, -17.96, -18.28, -18.675, -19.345, -19.56, -19.125, -19.805, 
    -19.305, -14.49, -11.81, -11.34, -11.38, -10.775, -10.575, -10.95, 
    -12.405, -14.26, -15.32, -16.83, -15.885, -16.525, -16.755, -16.51, 
    -15.7, -15.335, -15.35, -15.14, -14.785, -14.17, -13.585, -13.835, 
    -14.24, -12.725, -10.805, -9.535, -7.9, -7.18, -6.33, -7.795, -9.215, 
    -10.115, -9.975, -9.47, -9.36, -9.225, -8.995, -9.485, -9.485, -9.63, 
    -10.185, -11.245, -9.905, -9.77, -10.84, -12.165, -12.645, -12.71, 
    -12.485, -11.98, -10.905, -10.755, -11.565, -12.84, -14.165, -15.435, 
    -15.755, -15.655, -16.355, -17.17, -16.77, -16.02, -15.865, -16.38, 
    -17.825, -18.595, -19.02, -19.315, -19.555, -19.755, -19.985, -19.705, 
    -19.19, -18.81, -18.725, -18.26, -18.495, -18.97, -19.66, -20.705, 
    -21.335, -21.745, -22.295, -23.25, -24.245, -24.665, -24.505, -24.485, 
    -24.37, -24.205, -23.345, -22.25, -22.24, -22.17, -22.07, -21.72, 
    -18.895, -19.35, -17.555, -14.885, -12.675, -15.025, -18.625, -17.785, 
    -16.245, -17.095, -16.09, -16.875, -17.51, -18.045, -18.28, -18.3, 
    -18.415, -17.535, -16.975, -17.025, -17.1, -17.755, -18.285, -18.105, 
    -18.125, -17.525, -17.12, -17.48, -18.1, -18.54, -19.775, -20.585, 
    -21.17, -21.385, -21.095, -21.08, -21.235, -20.99, -20.805, -20.515, 
    -20.42, -20.185, -20.075, -20.405, -20.71, -21.015, -20.97, -20.575, 
    -20.225, -19.76, -19.475, -19.22, -19.465, -19.27, -19.115, -19.405, 
    -19.44, -19.37, -19.37, -19.395, -19.415, -19.415, -19.275, -19.17, 
    -19.21, -19.08, -18.99, -18.95, -18.815, -19.28, -18.905, -15.135, 
    -12.275, -11.595, -10.325, -10.455, -11.855, -12.435, -14.485, -15.87, 
    -17.055, -16.975, -16.375, -16.115, -16.07, -16, -15.48, -15.11, -14.535, 
    -14.875, -14.745, -14.215, -13.755, -13.425, -12.825, -10.51, -7.39, 
    -5.575, -4.445, -4.69, -4.975, -6.65, -7.895, -9.725, -11.065, -10.655, 
    -11.37, -10.1, -9.975, -9.885, -9.42, -9.41, -8.945, -8.61, -8.47, 
    -8.175, -7.835, -7.43, -7.385, -7.315, -6.92, -6.52, -6.23, -5.77, -5.79, 
    -6.225, -6.285, -6.125, -5.98, -5.755, -5.645, -5.51, -5.42, -5.425, 
    -5.535, -5.615, -5.5, -5.315, -5.195, -5.08, -5.12, -5.225, -5.365, 
    -5.59, -5.365, -5.44, -5.41, -5.505, -5.91, -6.135, -6.27, -6.38, -6.515, 
    -6.58, -6.55, -6.56, -6.645, -6.965, -7.265, -7.38, -7.825, -7.89, -7.78, 
    -7.7, -7.755, -7.95, -8.075, -8.12, -8.325, -8.255, -7.81, -8.43, -8.73, 
    -8.65, -9.255, -9.505, -9.465, -9.515, -9.92, -10.06, -10.07, -10.025, 
    -9.935, -9.81, -9.62, -8.785, -8.325, -8.485, -8.735, -8.785, -8.92, 
    -5.815, -4.445, -2.155, -2.13, -4.205, -4.08, -5.545, -6.225, -6.72, 
    -6.51, -6.09, -5.84, -5.775, -5.79, -5.185, -5.145, -4.935, -4.48, -4.06, 
    -3.765, -3.84, -4.545, -4.635, -3.765, -2.795, -2.095, -2.21, -2.855, 
    -3.545, -3.3, -3.06, -2.925, -3.525, -3.695, -3.95, -3.685, -3.495, 
    -3.18, -2.925, -3.41, -3.555, -3.325, -3.215, -3.42, -3.67, -3.945, 
    -4.09, -4.305, -4.125, -3.16, -3.65, -3.36, -2.73, -2.61, -3.21, -4.645, 
    -5.35, -5.675, -5.55, -5.51, -5.575, -5.635, -6.055, -6.94, -7.69, 
    -8.405, -9.185, -8.205, -7.705, -7.895, -7.725, -7.58, -6.49, -3.005, 
    -4.335, -3.93, -4.2, -3.965, -5.115, -6.095, -7.21, -7.88, -8.145, 
    -8.285, -8.885, -8.875, -8.96, -9.115, -8.93, -9.305, -9.47, -9.33, 
    -7.835, -7.315, -7.565, -7.18, -6.55, -5.3, -4.76, -4.48, -4.66, -4.61, 
    -4.58, -4.835, -5.255, -5.445, -5.325, -5.35, -5.245, -5.005, -4.79, 
    -4.74, -4.655, -4.06, -3.845, -3.125, -3.29, -2.995, -3.185, -3.31, 
    -2.025, 1.175, 2.505, 3.175, 3.145, 2.57, 1.095, -1.35, -2.875, -3.63, 
    -4.415, -5.305, -5.74, -4.94, -4.63, -4.425, -4.875, -5.035, -4.79, 
    -5.865, -5.805, -5.955, -5.34, -5.38, -2.91, -0.385, -0.27, 0.215, -0.42, 
    -0.215, -1.255, -2.87, -4.465, -5.465, -7.125, -7.495, -6.945, -5.57, 
    -5.24, -4.35, -4.25, -4.575, -4.62, -4.525, -4.58, -5.09, -5.075, -5.31, 
    -5.065, -4.22, -4.815, -5.265, -5.525, -6.25, -6.02, -6.115, -6.55, 
    -6.92, -6.215, -5.89, -5.82, -5.755, -5.795, -6.735, -8.43, -9.43, -8.76, 
    -8.13, -7.59, -7.745, -8.195, -8.035, -7.89, -7.93, -8.515, -8.45, -8.89, 
    -9.35, -10.29, -11.62, -12.92, -13.94, -14.675, -15.21, -16, -16.61, 
    -16.38, -17.19, -17.32, -17.855, -17.57, -18.915, -18.505, -17.815, 
    -18.93, -19.07, -15.53, -13.015, -12.67, -12.56, -12.655, -11.455, 
    -12.965, -14.29, -15.45, -15.815, -15.785, -15.355, -14.63, -14.145, 
    -14.09, -14.285, -14.1, -13.745, -13.875, -14.36, -14.435, -13.25, -12.4, 
    -12.58, -11.29, -8.965, -8.625, -8.975, -9.55, -10.125, -11.08, -11.315, 
    -12.695, -13.315, -13.875, -13.795, -14.37, -14.84, -13.87, -13.465, 
    -13.915, -14.755, -15.205, -15.305, -15.57, -15.355, -15.43, -14.65, 
    -9.12, -4.545, -3, -5.655, -6.365, -6.82, -6.97, -8.125, -10.44, -12.505, 
    -12.785, -12.57, -11.98, -11.945, -12.24, -11.8, -11.285, -10.035, 
    -10.09, -9.615, -10.11, -10.335, -9.92, -10.165, -7.91, -5.725, -5.41, 
    -5.31, -5.18, -5.97, -6.53, -7.595, -8.935, -9.815, -10.375, -10.545, 
    -11.495, -11.895, -12.705, -12.995, -12.85, -13.365, -12.865, -13.145, 
    -13.335, -13.625, -11.99, -12.155, -7.805, -2.85, -2.62, -2.51, -2.495, 
    -2.89, -3.86, -5.75, -8.58, -10.49, -9.89, -9.2, -9.57, -9.025, -9.41, 
    -9.21, -10.37, -10.85, -10.56, -9.405, -9.39, -10.125, -10.545, -9.535, 
    -8.555, -7.765, -8.935, -8.975, -8.225, -8.225, -8.305, -9.36, -10.3, 
    -10.46, -10.32, -10.325, -10.44, -10.57, -10.73, -10.81, -10.83, -10.85, 
    -10.68, -10.515, -10.485, -10.46, -10.375, -10.2, -9.87, -9.71, -9.97, 
    -10.115, -10.29, -10.265, -10.525, -10.655, -10.83, -11.13, -11.32, 
    -11.45, -11.365, -11.41, -11.175, -11, -11.05, -11.16, -11.21, -11.25, 
    -11.325, -11.46, -11.74, -11.78, -11.23, -10.245, -9.775, -9.115, -8.925, 
    -10.265, -10.64, -11.025, -11.22, -11.205, -11.165, -11, -10.64, -10.21, 
    -9.67, -8.725, -7.44, -7.26, -7.165, -6.45, -6.07, -5.98, -5.965, -5.635, 
    -4.63, -3.835, -3.85, -3.82, -4.06, -3.585, -4.02, -4.765, -5.095, -5.26, 
    -5.36, -5, -4.545, -4.355, -4.075, -4.35, -4.48, -4.435, -4.39, -4.57, 
    -4.73, -5.175, -5.51, -6.235, -6.595, -6.35, -6.12, -6.375, -5.735, 
    -6.26, -6.19, -6.82, -7.175, -7.385, -7.775, -8.295, -8.16, -8.425, 
    -8.16, -7.82, -7.76, -7.835, -7.975, -8.065, -8.135, -8.09, -7.875, 
    -7.91, -7.56, -6.925, -5.675, -5.265, -4.71, -4.275, -5.165, -7.075, 
    -7.53, -8.385, -10.07, -11.04, -9.97, -9.465, -9.525, -9.72, -9.175, 
    -8.805, -9.18, -8.68, -9.065, -9.46, -9.745, -8.465, -6.73, -3.945, 
    -0.485, -0.495, -0.645, -2.17, -4.61, -5.76, -6.04, -6.25, -6.28, -5.96, 
    -6.185, -5.615, -5.485, -5.62, -5.33, -5.25, -5.07, -4.695, -4.665, 
    -4.62, -4.345, -4.385, -4.2, -4.09, -4.535, -3.27, -3.08, -3.26, -3.99, 
    -4.615, -5.075, -5.045, -4.375, -4.35, -4.355, -4.49, -4.785, -4.645, 
    -4.725, -4.53, -4.265, -4.075, -3.99, -3.95, -3.695, -3.64, -3.775, 
    -3.84, -3.81, -3.76, -3.865, -4.39, -4.74, -5.52, -6.44, -7.42, -7.99, 
    -8.725, -10.68, -12.035, -12.77, -12.49, -13.635, -15.155, -15.77, 
    -16.06, -16.15, -15.66, -15.92, -15.74, -12.88, -9.905, -6.055, -4.78, 
    -5.285, -5.765, -7.07, -8.32, -10.375, -12.445, -12.86, -12.95, -13.015, 
    -12.6, -12.31, -11.595, -11.38, -11.495, -11.11, -11.01, -10.505, -10.46, 
    -10.64, -10.375, -7.355, -3.06, -0.025, 0.585, -1.085, -1.615, -2.14, 
    -2.935, -4.09, -4.345, -5.01, -4.615, -4.715, -4.73, -4.525, -4.585, 
    -4.71, -5.085, -4.83, -4.06, -4.135, -4.375, -4.645, -5.415, -4.645, 
    -2.545, -1.125, -0.895, -0.94, -1.635, -2.395, -2.705, -3.54, -4.98, 
    -4.475, -4.38, -4.09, -5.535, -5.845, -5.85, -4.81, -4.02, -4.13, -4.63, 
    -5.645, -5.195, -5.64, -5.865, -2.765, 0.66, 1.53, 1.22, 1.9, 1.68, 1.07, 
    -0.37, -1.655, -3.4, -4.36, -4.665, -4.765, -4.8, -4.94, -5.55, -5.315, 
    -5.13, -4.915, -5.165, -5.695, -5.65, -5.645, -5.63, -1.34, 2.43, 3.78, 
    4.19, 3.38, 3.8, 3.395, 1.47, 0.345, -0.085, -0.675, -0.12, -2.305, 
    -4.25, -4.78, -4.225, -4.34, -5.215, -5.575, -2.12, -3.445, -1.35, 
    -0.435, -0.095, 1.43, 1.76, 2.09, 2.54, 2.19, 1.905, 1.185, 1.175, 
    -0.655, -1.435, -2.045, -1.88, -3.135, -3.9, -3.785, -2.76, -2.755, 
    -2.575, -3.11, -4.3, -5.945, -6.455, -6.14, -5.77, -3.155, 0.405, 2.715, 
    2.23, 2.61, 0.42, 1.26, -0.115, -1.685, -2.155, -2.805, -3.24, -3.125, 
    -3.45, -4.3, -4.965, -5.03, -5.665, -5.7, -5.585, -5.795, -5.925, -6.055, 
    -6.155, -5.78, -5.09, -5.12, -4.5, -4.32, -4.195, -4.57, -5.32, -6.03, 
    -6.63, -7.41, -8.055, -8.335, -8.65, -8.58, -8.6, -9.29, -10.37, -10.12, 
    -9.49, -8.435, -8.325, -9.545, -7.535, -6.17, -4.84, -3.28, -2.545, 
    -2.07, -1.18, -1.835, -2.55, -2.56, -2.47, -2.72, -2.68, -3.175, -3.03, 
    -2.35, -2.535, -3.365, -3.07, -3.2, -3.105, -4.345, -3.715, -3.79, 
    -3.585, -1.015, 0.52, 2.87, 3.41, 2.845, 1.565, 1.67, 0.03, -2.025, 
    -2.87, -3.785, -3.61, -3.735, -3.275, -2.905, -3.425, -2.73, -3.705, 
    -3.81, -4.375, -5.085, -6.665, -5.465, -4.25, -1.75, 1.065, 0.805, 1.4, 
    2.235, 2.115, 1.685, -0.19, -2.595, -4.095, -4.015, -3.665, -3.205, 
    -3.03, -2.985, -3.485, -4.155, -4.565, -5.53, -5.695, -4.95, -5.59, 
    -5.92, -5.84, -5.445, -4.705, -4.615, -3.24, -3.86, -3.725, -4.13, -4.04, 
    -4.295, -4.435, -4.19, -4.33, -4.815, -5.005, -5.065, -4.825, -4.8, 
    -4.64, -4.24, -4.485, -4.825, -4.995, -5.245, -5.265, -5.22, -5.775, 
    -5.79, -5.325, -4.55, -5.65, -5.77, -5.91, -7.145, -7.855, -9.365, -8.31, 
    -7.795, -7.275, -7.145, -7.52, -7.775, -7.36, -7.85, -8.25, -8.15, -8.14, 
    -8.6, -8.595, -7.36, -5.85, -4.705, -5.065, -5.045, -5.975, -5.795, 
    -5.55, -6.68, -7.605, -8.11, -7.86, -7.685, -7.485, -7.135, -7.315, 
    -7.36, -7.205, -6.965, -6.82, -6.835, -6.99, -6.895, -6.84, -6.525, 
    -6.02, -5.675, -4.24, -4.675, -4.665, -4.695, -5.27, -6.405, -7.235, 
    -7.1, -7.345, -7.725, -7.48, -7.275, -7.79, -7.68, -7.6, -7.385, -6.56, 
    -5.955, -6.11, -6.545, -6.635, -6.515, -6.17, -5.305, -5.655, -6.005, 
    -6.695, -7.035, -7.16, -7.205, -7.37, -7.59, -7.7, -7.82, -8.26, -8.495, 
    -8.565, -8.605, -8.81, -9.19, -9.41, -9.475, -9.51, -9.555, -9.64, -9.5, 
    -9.35, -9.2, -9.22, -9.44, -9.615, -9.78, -9.78, -9.685, -9.65, -9.625, 
    -9.6, -9.625, -9.74, -9.875, -9.965, -10.075, -10.175, -10.23, -10.215, 
    -10.255, -10.31, -10.31, -10.375, -10.22, -9.755, -8.63, -7.215, -8.505, 
    -9.28, -9.46, -10.105, -10.5, -10.91, -11.29, -11.585, -11.655, -11.925, 
    -12.14, -12.165, -11.54, -11.055, -11.17, -11.26, -10.815, -10.49, 
    -10.505, -10.025, -9.39, -9.115, -8.83, -8.345, -6.725, -6.045, -5.165, 
    -5.88, -7.2, -7.63, -7.795, -8.485, -10.6, -11.19, -9.17, -8.75, -9.605, 
    -10.255, -10.735, -10.06, -8.325, -6.455, -6.355, -6.43, -5.34, -3.955, 
    -2.875, -3.755, -3.085, -2.67, -2.3, -3.165, -4.445, -5.105, -5.345, 
    -5.525, -6.06, -6.5, -7.16, -7.35, -7.11, -8.16, -8.68, -8.495, -8.6, 
    -8.165, -7.945, -8.435, -6.715, -4.175, -2.98, -2.245, -2.635, -2.99, 
    -3.59, -4.015, -5.26, -6.64, -6.955, -6.945, -6.925, -6.8, -7.245, -7.65, 
    -8, -8.105, -8.07, -7.99, -8.055, -8.935, -9.44, -9.425, -6.345, -4.485, 
    -3.795, -3.12, -2.88, -2.25, -2.125, -3.3, -5.79, -7.66, -8.255, -8.985, 
    -9.48, -9.625, -10.43, -10.325, -9.5, -10.63, -10.7, -10.325, -10.52, 
    -10.815, -10.675, -10.165, -6.18, -3.14, -1.37, -1.145, -0.9, -0.62, 
    -0.66, -3.105, -4.88, -6.73, -6.945, -7.765, -8.805, -8.975, -8.825, 
    -8.2, -7.88, -9.39, -8.385, -8.9, -7.305, -7.37, -9.75, -9.985, -6.56, 
    -1.025, 1.22, 1.44, 0.785, 0.615, 0.5, -1.65, -3.605, -4.805, -5.71, 
    -5.435, -5.24, -5.53, -5.61, -5.725, -6.06, -6.46, -6.985, -7.275, 
    -7.265, -7.285, -7.25, -7.255, -7.085, -6.685, -6.695, -6.635, -6.77, 
    -6.92, -6.815, -7.225, -7.32, -7.365, -7.32, -7.345, -7.475, -7.72, 
    -7.725, -7.9, -8.01, -8.005, -8.005, -8.155, -8.295, -8.405, -8.615, 
    -8.675, -8.375, -7.33, -6.57, -6.145, -7.515, -6.66, -5.42, -6.335, 
    -7.645, -8.825, -9.915, -11.955, -11.91, -11.31, -10.255, -10.925, 
    -10.965, -10.295, -9.375, -9.245, -9.375, -9.755, -10.95, -10.68, -6.425, 
    -0.755, -0.125, -1.15, -2.785, -3.34, -3.385, -3.89, -4.725, -6.705, 
    -7.995, -7.465, -7.3, -7.64, -9.24, -9.84, -10.31, -9.99, -9.83, -9.6, 
    -9.3, -8.495, -7.625, -6.185, -4.885, -5.4, -4.21, -1.24, -1.065, -1.255, 
    -1.425, -2.215, -3.815, -5.24, -5.98, -5.975, -6.325, -6.35, -6.46, 
    -6.48, -6.93, -7.535, -7.795, -8.035, -8.045, -7.93, -8.735, -8.93, 
    -7.295, -6.155, -6.31, -5.095, -4.445, -5.165, -6.095, -5.32, -6.735, 
    -8.38, -9.31, -9.57, -9.25, -9.895, -9.365, -8.545, -8.21, -7.295, -6.67, 
    -7.195, -6.61, -6.67, -6.725, -6.145, -5.555, -5.355, -4.36, -3.695, 
    -4.14, -4.485, -4.5, -4.57, -4.555, -4.615, -4.52, -4.37, -4.4, -4.33, 
    -4.315, -4.195, -4.16, -4.23, -4.41, -4.47, -4.605, -4.95, -5.225, -4.84, 
    -4, -3.795, -2.98, -1.985, -2.375, -2.63, -2.42, -2.535, -4.08, -6.485, 
    -6.71, -5.935, -6.07, -6.475, -6.465, -6.67, -6.925, -7.095, -7.7, -7.6, 
    -7.435, -7.48, -7.89, -8.11, -8.09, -8, -7.58, -7.225, -6.825, -6.825, 
    -6.71, -6.68, -7.045, -8.085, -8.965, -9.575, -9.685, -9.85, -10.19, 
    -10.47, -11.075, -11.385, -11.22, -12.165, -12.885, -14.19, -14.465, 
    -13.165, -6.15, -5.99, -6.675, -5.78, -4.725, -6.39, -7.43, -8.135, 
    -8.98, -10.35, -10.75, -11.035, -12.695, -13.41, -13.825, -14.255, 
    -14.295, -14.6, -15.105, -13.685, -12.32, -11.06, -11.32, -10.655, -9.62, 
    -9.305, -8.37, -8.195, -6.635, -8.045, -7.84, -7.43, -8.675, -11.25, 
    -13.195, -11.835, -12.225, -12.505, -11.32, -11.215, -10.7, -10.465, 
    -10.26, -9.855, -9.795, -9.725, -9.865, -9.715, -8.72, -8.1, -7.4, -6.72, 
    -6.94, -8.03, -7.95, -7.94, -8.505, -8.735, -8.84, -8.865, -9.165, -9.31, 
    -9.26, -9.06, -9.1, -9.045, -8.615, -8.56, -8.64, -8.805, -8.88, -8.76, 
    -8.4, -7.845, -7.49, -7.125, -7.01, -6.955, -6.95, -6.745, -6.995, -7.18, 
    -7.28, -7.07, -7.095, -7.025, -6.625, -6.395, -6.305, -6.3, -6.215, 
    -6.22, -6.33, -6.355, -6.22, -5.985, -5.475, -5.3, -5.195, -4.985, -4.92, 
    -4.855, -5.115, -5.4, -5.455, -5.76, -5.695, -5.47, -5.305, -5.165, 
    -5.085, -5.23, -5.325, -5.285, -5.295, -5.315, -5.375, -5.275, -5.255, 
    -5.175, -4.885, -4.745, -4.825, -4.745, -4.745, -4.535, -5.295, -5.79, 
    -6.865, -8.16, -8.745, -9.715, -10.79, -9.655, -10.88 ;
}
